module main (
    input wire clock,
    input wire reset,
    input wire [7:0] a,
    input wire [7:0] b,
    input wire [7:0] c,
    input wire [7:0] d,
    input wire [7:0] e,
    input wire [7:0] f,
    input wire [7:0] g,
    input wire [7:0] h,
    input wire en,
    output wire [7:0] y
);
    wire gnd;
    wire vcc;
    wire t2;
    wire t3;
    wire t4;
    wire t5;
    wire t6;
    wire t7;
    wire t8;
    wire t9;
    wire t10;
    wire t11;
    wire t12;
    wire t13;
    wire t14;
    wire t15;
    wire t16;
    wire t17;
    wire t18;
    wire t19;
    wire t20;
    wire t21;
    wire t22;
    wire t23;
    wire t24;
    wire t25;
    wire [7:0] t26;
    wire [7:0] t27;
    wire t28;
    wire t29;
    wire t30;
    wire t31;
    wire t32;
    wire t33;
    wire t34;
    wire t35;
    wire t36;
    wire t37;
    wire t38;
    wire t39;
    wire t40;
    wire t41;
    wire t42;
    wire t43;
    wire t46;
    wire t47;
    wire t48;
    wire t49;
    wire t50;
    wire t51;
    wire t52;
    wire t53;
    wire t54;
    wire t55;
    wire t56;
    wire t57;
    wire t58;
    wire t59;
    wire t60;
    wire t61;
    wire t62;
    wire t63;
    wire t64;
    wire t65;
    wire t66;
    wire t67;
    wire t68;
    wire t69;
    wire [7:0] t70;
    wire [7:0] t71;
    wire t72;
    wire t73;
    wire t74;
    wire t75;
    wire t76;
    wire t77;
    wire t78;
    wire t79;
    wire t80;
    wire t81;
    wire t82;
    wire t83;
    wire t84;
    wire t85;
    wire t86;
    wire t87;
    wire [7:0] t0;
    wire t90;
    wire t91;
    wire t92;
    wire t93;
    wire t94;
    wire t95;
    wire t96;
    wire t97;
    wire t98;
    wire t99;
    wire t100;
    wire t101;
    wire t102;
    wire t103;
    wire t104;
    wire t105;
    wire t106;
    wire t107;
    wire t108;
    wire t109;
    wire t110;
    wire t111;
    wire t112;
    wire t113;
    wire [7:0] t114;
    wire [7:0] t115;
    wire t116;
    wire t117;
    wire t118;
    wire t119;
    wire t120;
    wire t121;
    wire t122;
    wire t123;
    wire t124;
    wire t125;
    wire t126;
    wire t127;
    wire t128;
    wire t129;
    wire t130;
    wire t131;
    wire [7:0] t1;
    wire t132;
    wire t133;
    wire t134;
    wire t135;
    wire t136;
    wire t137;
    wire t138;
    wire t139;
    wire t140;
    wire t141;
    wire t142;
    wire t143;
    wire t144;
    wire t145;
    wire t146;
    wire t147;
    wire t148;
    wire t149;
    wire t150;
    wire t151;
    wire t152;
    wire t153;
    wire t154;
    wire t155;
    wire [7:0] t156;
    wire [7:0] t157;
    wire t158;
    wire t159;
    wire t160;
    wire t161;
    wire t162;
    wire t163;
    wire t164;
    wire t165;
    wire t166;
    wire t167;
    wire t168;
    wire t169;
    wire t170;
    wire t171;
    wire t172;
    wire t173;
    wire [7:0] t44;
    wire t174;
    wire t175;
    wire t176;
    wire t177;
    wire t178;
    wire t179;
    wire t180;
    wire t181;
    wire t182;
    wire t183;
    wire t184;
    wire t185;
    wire t186;
    wire t187;
    wire t188;
    wire t189;
    wire t190;
    wire t191;
    wire t192;
    wire t193;
    wire t194;
    wire t195;
    wire t196;
    wire t197;
    wire [7:0] t198;
    wire [7:0] t199;
    wire t200;
    wire t201;
    wire t202;
    wire t203;
    wire t204;
    wire t205;
    wire t206;
    wire t207;
    wire t208;
    wire t209;
    wire t210;
    wire t211;
    wire t212;
    wire t213;
    wire t214;
    wire t215;
    wire [7:0] t45;
    wire t216;
    wire t217;
    wire t218;
    wire t219;
    wire t220;
    wire t221;
    wire t222;
    wire t223;
    wire t224;
    wire t225;
    wire t226;
    wire t227;
    wire t228;
    wire t229;
    wire t230;
    wire t231;
    wire t232;
    wire t233;
    wire t234;
    wire t235;
    wire t236;
    wire t237;
    wire t238;
    wire t239;
    wire [7:0] t240;
    wire [7:0] t241;
    wire t242;
    wire t243;
    wire t244;
    wire t245;
    wire t246;
    wire t247;
    wire t248;
    wire t249;
    wire t250;
    wire t251;
    wire t252;
    wire t253;
    wire t254;
    wire t255;
    wire t256;
    wire t257;
    wire [7:0] t88;
    wire t258;
    wire t259;
    wire t260;
    wire t261;
    wire t262;
    wire t263;
    wire t264;
    wire t265;
    wire t266;
    wire t267;
    wire t268;
    wire t269;
    wire t270;
    wire t271;
    wire t272;
    wire t273;
    wire t274;
    wire t275;
    wire t276;
    wire t277;
    wire t278;
    wire t279;
    wire t280;
    wire t281;
    wire [7:0] t282;
    wire [7:0] t283;
    wire t284;
    wire t285;
    wire t286;
    wire t287;
    wire t288;
    wire t289;
    wire t290;
    wire t291;
    wire t292;
    wire t293;
    wire t294;
    wire t295;
    wire t296;
    wire t297;
    wire t298;
    wire t299;
    wire [7:0] t89;
    GND _gnd (
        .G(gnd)
    );
    VCC _vcc (
        .P(vcc)
    );
    assign t2 = t0[0];
    assign t3 = t0[1];
    assign t4 = t0[2];
    assign t5 = t0[3];
    assign t6 = t0[4];
    assign t7 = t0[5];
    assign t8 = t0[6];
    assign t9 = t0[7];
    assign t10 = t1[0];
    assign t11 = t1[1];
    assign t12 = t1[2];
    assign t13 = t1[3];
    assign t14 = t1[4];
    assign t15 = t1[5];
    assign t16 = t1[6];
    assign t17 = t1[7];
    (*LOC = "SLICE_X0Y0", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t18 (
        .I0(t2),
        .I1(t10),
        .O(t18)
    );
    (*LOC = "SLICE_X0Y0", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t19 (
        .I0(t3),
        .I1(t11),
        .O(t19)
    );
    (*LOC = "SLICE_X0Y0", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t20 (
        .I0(t4),
        .I1(t12),
        .O(t20)
    );
    (*LOC = "SLICE_X0Y0", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t21 (
        .I0(t5),
        .I1(t13),
        .O(t21)
    );
    (*LOC = "SLICE_X0Y0", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t22 (
        .I0(t6),
        .I1(t14),
        .O(t22)
    );
    (*LOC = "SLICE_X0Y0", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t23 (
        .I0(t7),
        .I1(t15),
        .O(t23)
    );
    (*LOC = "SLICE_X0Y0", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t24 (
        .I0(t8),
        .I1(t16),
        .O(t24)
    );
    (*LOC = "SLICE_X0Y0", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t25 (
        .I0(t9),
        .I1(t17),
        .O(t25)
    );
    assign t26 = {t25, t24, t23, t22, t21, t20, t19, t18};
    (*LOC = "SLICE_X0Y0", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t27 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(t0),
        .O(t27),
        .S(t26)
    );
    assign t28 = t27[0];
    assign t29 = t27[1];
    assign t30 = t27[2];
    assign t31 = t27[3];
    assign t32 = t27[4];
    assign t33 = t27[5];
    assign t34 = t27[6];
    assign t35 = t27[7];
    (*LOC = "SLICE_X0Y0", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t36 (
        .C(clock),
        .CE(en),
        .D(t28),
        .Q(t36),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t37 (
        .C(clock),
        .CE(en),
        .D(t29),
        .Q(t37),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t38 (
        .C(clock),
        .CE(en),
        .D(t30),
        .Q(t38),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t39 (
        .C(clock),
        .CE(en),
        .D(t31),
        .Q(t39),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t40 (
        .C(clock),
        .CE(en),
        .D(t32),
        .Q(t40),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t41 (
        .C(clock),
        .CE(en),
        .D(t33),
        .Q(t41),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t42 (
        .C(clock),
        .CE(en),
        .D(t34),
        .Q(t42),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y0", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t43 (
        .C(clock),
        .CE(en),
        .D(t35),
        .Q(t43),
        .R(reset)
    );
    assign y = {t43, t42, t41, t40, t39, t38, t37, t36};
    assign t46 = t44[0];
    assign t47 = t44[1];
    assign t48 = t44[2];
    assign t49 = t44[3];
    assign t50 = t44[4];
    assign t51 = t44[5];
    assign t52 = t44[6];
    assign t53 = t44[7];
    assign t54 = t45[0];
    assign t55 = t45[1];
    assign t56 = t45[2];
    assign t57 = t45[3];
    assign t58 = t45[4];
    assign t59 = t45[5];
    assign t60 = t45[6];
    assign t61 = t45[7];
    (*LOC = "SLICE_X0Y1", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t62 (
        .I0(t46),
        .I1(t54),
        .O(t62)
    );
    (*LOC = "SLICE_X0Y1", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t63 (
        .I0(t47),
        .I1(t55),
        .O(t63)
    );
    (*LOC = "SLICE_X0Y1", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t64 (
        .I0(t48),
        .I1(t56),
        .O(t64)
    );
    (*LOC = "SLICE_X0Y1", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t65 (
        .I0(t49),
        .I1(t57),
        .O(t65)
    );
    (*LOC = "SLICE_X0Y1", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t66 (
        .I0(t50),
        .I1(t58),
        .O(t66)
    );
    (*LOC = "SLICE_X0Y1", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t67 (
        .I0(t51),
        .I1(t59),
        .O(t67)
    );
    (*LOC = "SLICE_X0Y1", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t68 (
        .I0(t52),
        .I1(t60),
        .O(t68)
    );
    (*LOC = "SLICE_X0Y1", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t69 (
        .I0(t53),
        .I1(t61),
        .O(t69)
    );
    assign t70 = {t69, t68, t67, t66, t65, t64, t63, t62};
    (*LOC = "SLICE_X0Y1", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t71 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(t44),
        .O(t71),
        .S(t70)
    );
    assign t72 = t71[0];
    assign t73 = t71[1];
    assign t74 = t71[2];
    assign t75 = t71[3];
    assign t76 = t71[4];
    assign t77 = t71[5];
    assign t78 = t71[6];
    assign t79 = t71[7];
    (*LOC = "SLICE_X0Y1", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t80 (
        .C(clock),
        .CE(en),
        .D(t72),
        .Q(t80),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t81 (
        .C(clock),
        .CE(en),
        .D(t73),
        .Q(t81),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t82 (
        .C(clock),
        .CE(en),
        .D(t74),
        .Q(t82),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t83 (
        .C(clock),
        .CE(en),
        .D(t75),
        .Q(t83),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t84 (
        .C(clock),
        .CE(en),
        .D(t76),
        .Q(t84),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t85 (
        .C(clock),
        .CE(en),
        .D(t77),
        .Q(t85),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t86 (
        .C(clock),
        .CE(en),
        .D(t78),
        .Q(t86),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y1", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t87 (
        .C(clock),
        .CE(en),
        .D(t79),
        .Q(t87),
        .R(reset)
    );
    assign t0 = {t87, t86, t85, t84, t83, t82, t81, t80};
    assign t90 = t88[0];
    assign t91 = t88[1];
    assign t92 = t88[2];
    assign t93 = t88[3];
    assign t94 = t88[4];
    assign t95 = t88[5];
    assign t96 = t88[6];
    assign t97 = t88[7];
    assign t98 = t89[0];
    assign t99 = t89[1];
    assign t100 = t89[2];
    assign t101 = t89[3];
    assign t102 = t89[4];
    assign t103 = t89[5];
    assign t104 = t89[6];
    assign t105 = t89[7];
    (*LOC = "SLICE_X0Y2", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t106 (
        .I0(t90),
        .I1(t98),
        .O(t106)
    );
    (*LOC = "SLICE_X0Y2", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t107 (
        .I0(t91),
        .I1(t99),
        .O(t107)
    );
    (*LOC = "SLICE_X0Y2", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t108 (
        .I0(t92),
        .I1(t100),
        .O(t108)
    );
    (*LOC = "SLICE_X0Y2", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t109 (
        .I0(t93),
        .I1(t101),
        .O(t109)
    );
    (*LOC = "SLICE_X0Y2", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t110 (
        .I0(t94),
        .I1(t102),
        .O(t110)
    );
    (*LOC = "SLICE_X0Y2", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t111 (
        .I0(t95),
        .I1(t103),
        .O(t111)
    );
    (*LOC = "SLICE_X0Y2", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t112 (
        .I0(t96),
        .I1(t104),
        .O(t112)
    );
    (*LOC = "SLICE_X0Y2", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t113 (
        .I0(t97),
        .I1(t105),
        .O(t113)
    );
    assign t114 = {t113, t112, t111, t110, t109, t108, t107, t106};
    (*LOC = "SLICE_X0Y2", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t115 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(t88),
        .O(t115),
        .S(t114)
    );
    assign t116 = t115[0];
    assign t117 = t115[1];
    assign t118 = t115[2];
    assign t119 = t115[3];
    assign t120 = t115[4];
    assign t121 = t115[5];
    assign t122 = t115[6];
    assign t123 = t115[7];
    (*LOC = "SLICE_X0Y2", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t124 (
        .C(clock),
        .CE(en),
        .D(t116),
        .Q(t124),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t125 (
        .C(clock),
        .CE(en),
        .D(t117),
        .Q(t125),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t126 (
        .C(clock),
        .CE(en),
        .D(t118),
        .Q(t126),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t127 (
        .C(clock),
        .CE(en),
        .D(t119),
        .Q(t127),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t128 (
        .C(clock),
        .CE(en),
        .D(t120),
        .Q(t128),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t129 (
        .C(clock),
        .CE(en),
        .D(t121),
        .Q(t129),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t130 (
        .C(clock),
        .CE(en),
        .D(t122),
        .Q(t130),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y2", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t131 (
        .C(clock),
        .CE(en),
        .D(t123),
        .Q(t131),
        .R(reset)
    );
    assign t1 = {t131, t130, t129, t128, t127, t126, t125, t124};
    assign t132 = a[0];
    assign t133 = a[1];
    assign t134 = a[2];
    assign t135 = a[3];
    assign t136 = a[4];
    assign t137 = a[5];
    assign t138 = a[6];
    assign t139 = a[7];
    assign t140 = b[0];
    assign t141 = b[1];
    assign t142 = b[2];
    assign t143 = b[3];
    assign t144 = b[4];
    assign t145 = b[5];
    assign t146 = b[6];
    assign t147 = b[7];
    (*LOC = "SLICE_X0Y3", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t148 (
        .I0(t132),
        .I1(t140),
        .O(t148)
    );
    (*LOC = "SLICE_X0Y3", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t149 (
        .I0(t133),
        .I1(t141),
        .O(t149)
    );
    (*LOC = "SLICE_X0Y3", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t150 (
        .I0(t134),
        .I1(t142),
        .O(t150)
    );
    (*LOC = "SLICE_X0Y3", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t151 (
        .I0(t135),
        .I1(t143),
        .O(t151)
    );
    (*LOC = "SLICE_X0Y3", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t152 (
        .I0(t136),
        .I1(t144),
        .O(t152)
    );
    (*LOC = "SLICE_X0Y3", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t153 (
        .I0(t137),
        .I1(t145),
        .O(t153)
    );
    (*LOC = "SLICE_X0Y3", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t154 (
        .I0(t138),
        .I1(t146),
        .O(t154)
    );
    (*LOC = "SLICE_X0Y3", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t155 (
        .I0(t139),
        .I1(t147),
        .O(t155)
    );
    assign t156 = {t155, t154, t153, t152, t151, t150, t149, t148};
    (*LOC = "SLICE_X0Y3", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t157 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(a),
        .O(t157),
        .S(t156)
    );
    assign t158 = t157[0];
    assign t159 = t157[1];
    assign t160 = t157[2];
    assign t161 = t157[3];
    assign t162 = t157[4];
    assign t163 = t157[5];
    assign t164 = t157[6];
    assign t165 = t157[7];
    (*LOC = "SLICE_X0Y3", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t166 (
        .C(clock),
        .CE(en),
        .D(t158),
        .Q(t166),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t167 (
        .C(clock),
        .CE(en),
        .D(t159),
        .Q(t167),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t168 (
        .C(clock),
        .CE(en),
        .D(t160),
        .Q(t168),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t169 (
        .C(clock),
        .CE(en),
        .D(t161),
        .Q(t169),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t170 (
        .C(clock),
        .CE(en),
        .D(t162),
        .Q(t170),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t171 (
        .C(clock),
        .CE(en),
        .D(t163),
        .Q(t171),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t172 (
        .C(clock),
        .CE(en),
        .D(t164),
        .Q(t172),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y3", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t173 (
        .C(clock),
        .CE(en),
        .D(t165),
        .Q(t173),
        .R(reset)
    );
    assign t44 = {t173, t172, t171, t170, t169, t168, t167, t166};
    assign t174 = c[0];
    assign t175 = c[1];
    assign t176 = c[2];
    assign t177 = c[3];
    assign t178 = c[4];
    assign t179 = c[5];
    assign t180 = c[6];
    assign t181 = c[7];
    assign t182 = d[0];
    assign t183 = d[1];
    assign t184 = d[2];
    assign t185 = d[3];
    assign t186 = d[4];
    assign t187 = d[5];
    assign t188 = d[6];
    assign t189 = d[7];
    (*LOC = "SLICE_X0Y4", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t190 (
        .I0(t174),
        .I1(t182),
        .O(t190)
    );
    (*LOC = "SLICE_X0Y4", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t191 (
        .I0(t175),
        .I1(t183),
        .O(t191)
    );
    (*LOC = "SLICE_X0Y4", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t192 (
        .I0(t176),
        .I1(t184),
        .O(t192)
    );
    (*LOC = "SLICE_X0Y4", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t193 (
        .I0(t177),
        .I1(t185),
        .O(t193)
    );
    (*LOC = "SLICE_X0Y4", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t194 (
        .I0(t178),
        .I1(t186),
        .O(t194)
    );
    (*LOC = "SLICE_X0Y4", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t195 (
        .I0(t179),
        .I1(t187),
        .O(t195)
    );
    (*LOC = "SLICE_X0Y4", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t196 (
        .I0(t180),
        .I1(t188),
        .O(t196)
    );
    (*LOC = "SLICE_X0Y4", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t197 (
        .I0(t181),
        .I1(t189),
        .O(t197)
    );
    assign t198 = {t197, t196, t195, t194, t193, t192, t191, t190};
    (*LOC = "SLICE_X0Y4", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t199 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(c),
        .O(t199),
        .S(t198)
    );
    assign t200 = t199[0];
    assign t201 = t199[1];
    assign t202 = t199[2];
    assign t203 = t199[3];
    assign t204 = t199[4];
    assign t205 = t199[5];
    assign t206 = t199[6];
    assign t207 = t199[7];
    (*LOC = "SLICE_X0Y4", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t208 (
        .C(clock),
        .CE(en),
        .D(t200),
        .Q(t208),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t209 (
        .C(clock),
        .CE(en),
        .D(t201),
        .Q(t209),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t210 (
        .C(clock),
        .CE(en),
        .D(t202),
        .Q(t210),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t211 (
        .C(clock),
        .CE(en),
        .D(t203),
        .Q(t211),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t212 (
        .C(clock),
        .CE(en),
        .D(t204),
        .Q(t212),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t213 (
        .C(clock),
        .CE(en),
        .D(t205),
        .Q(t213),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t214 (
        .C(clock),
        .CE(en),
        .D(t206),
        .Q(t214),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y4", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t215 (
        .C(clock),
        .CE(en),
        .D(t207),
        .Q(t215),
        .R(reset)
    );
    assign t45 = {t215, t214, t213, t212, t211, t210, t209, t208};
    assign t216 = e[0];
    assign t217 = e[1];
    assign t218 = e[2];
    assign t219 = e[3];
    assign t220 = e[4];
    assign t221 = e[5];
    assign t222 = e[6];
    assign t223 = e[7];
    assign t224 = f[0];
    assign t225 = f[1];
    assign t226 = f[2];
    assign t227 = f[3];
    assign t228 = f[4];
    assign t229 = f[5];
    assign t230 = f[6];
    assign t231 = f[7];
    (*LOC = "SLICE_X0Y5", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t232 (
        .I0(t216),
        .I1(t224),
        .O(t232)
    );
    (*LOC = "SLICE_X0Y5", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t233 (
        .I0(t217),
        .I1(t225),
        .O(t233)
    );
    (*LOC = "SLICE_X0Y5", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t234 (
        .I0(t218),
        .I1(t226),
        .O(t234)
    );
    (*LOC = "SLICE_X0Y5", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t235 (
        .I0(t219),
        .I1(t227),
        .O(t235)
    );
    (*LOC = "SLICE_X0Y5", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t236 (
        .I0(t220),
        .I1(t228),
        .O(t236)
    );
    (*LOC = "SLICE_X0Y5", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t237 (
        .I0(t221),
        .I1(t229),
        .O(t237)
    );
    (*LOC = "SLICE_X0Y5", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t238 (
        .I0(t222),
        .I1(t230),
        .O(t238)
    );
    (*LOC = "SLICE_X0Y5", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t239 (
        .I0(t223),
        .I1(t231),
        .O(t239)
    );
    assign t240 = {t239, t238, t237, t236, t235, t234, t233, t232};
    (*LOC = "SLICE_X0Y5", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t241 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(e),
        .O(t241),
        .S(t240)
    );
    assign t242 = t241[0];
    assign t243 = t241[1];
    assign t244 = t241[2];
    assign t245 = t241[3];
    assign t246 = t241[4];
    assign t247 = t241[5];
    assign t248 = t241[6];
    assign t249 = t241[7];
    (*LOC = "SLICE_X0Y5", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t250 (
        .C(clock),
        .CE(en),
        .D(t242),
        .Q(t250),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t251 (
        .C(clock),
        .CE(en),
        .D(t243),
        .Q(t251),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t252 (
        .C(clock),
        .CE(en),
        .D(t244),
        .Q(t252),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t253 (
        .C(clock),
        .CE(en),
        .D(t245),
        .Q(t253),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t254 (
        .C(clock),
        .CE(en),
        .D(t246),
        .Q(t254),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t255 (
        .C(clock),
        .CE(en),
        .D(t247),
        .Q(t255),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t256 (
        .C(clock),
        .CE(en),
        .D(t248),
        .Q(t256),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y5", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t257 (
        .C(clock),
        .CE(en),
        .D(t249),
        .Q(t257),
        .R(reset)
    );
    assign t88 = {t257, t256, t255, t254, t253, t252, t251, t250};
    assign t258 = g[0];
    assign t259 = g[1];
    assign t260 = g[2];
    assign t261 = g[3];
    assign t262 = g[4];
    assign t263 = g[5];
    assign t264 = g[6];
    assign t265 = g[7];
    assign t266 = h[0];
    assign t267 = h[1];
    assign t268 = h[2];
    assign t269 = h[3];
    assign t270 = h[4];
    assign t271 = h[5];
    assign t272 = h[6];
    assign t273 = h[7];
    (*LOC = "SLICE_X0Y6", BEL = "A6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t274 (
        .I0(t258),
        .I1(t266),
        .O(t274)
    );
    (*LOC = "SLICE_X0Y6", BEL = "B6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t275 (
        .I0(t259),
        .I1(t267),
        .O(t275)
    );
    (*LOC = "SLICE_X0Y6", BEL = "C6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t276 (
        .I0(t260),
        .I1(t268),
        .O(t276)
    );
    (*LOC = "SLICE_X0Y6", BEL = "D6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t277 (
        .I0(t261),
        .I1(t269),
        .O(t277)
    );
    (*LOC = "SLICE_X0Y6", BEL = "E6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t278 (
        .I0(t262),
        .I1(t270),
        .O(t278)
    );
    (*LOC = "SLICE_X0Y6", BEL = "F6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t279 (
        .I0(t263),
        .I1(t271),
        .O(t279)
    );
    (*LOC = "SLICE_X0Y6", BEL = "G6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t280 (
        .I0(t264),
        .I1(t272),
        .O(t280)
    );
    (*LOC = "SLICE_X0Y6", BEL = "H6LUT"*)
    LUT2 # (
        .INIT(4'h6)
    ) __t281 (
        .I0(t265),
        .I1(t273),
        .O(t281)
    );
    assign t282 = {t281, t280, t279, t278, t277, t276, t275, t274};
    (*LOC = "SLICE_X0Y6", BEL = "CARRY8"*)
    CARRY8 # (
        .CARRY_TYPE("SINGLE_CY8")
    ) __t283 (
        .CI(1'b0),
        .CI_TOP(1'b0),
        .CO(),
        .DI(g),
        .O(t283),
        .S(t282)
    );
    assign t284 = t283[0];
    assign t285 = t283[1];
    assign t286 = t283[2];
    assign t287 = t283[3];
    assign t288 = t283[4];
    assign t289 = t283[5];
    assign t290 = t283[6];
    assign t291 = t283[7];
    (*LOC = "SLICE_X0Y6", BEL = "AFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t292 (
        .C(clock),
        .CE(en),
        .D(t284),
        .Q(t292),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "BFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t293 (
        .C(clock),
        .CE(en),
        .D(t285),
        .Q(t293),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "CFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t294 (
        .C(clock),
        .CE(en),
        .D(t286),
        .Q(t294),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "DFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t295 (
        .C(clock),
        .CE(en),
        .D(t287),
        .Q(t295),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "EFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t296 (
        .C(clock),
        .CE(en),
        .D(t288),
        .Q(t296),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "FFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t297 (
        .C(clock),
        .CE(en),
        .D(t289),
        .Q(t297),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "GFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t298 (
        .C(clock),
        .CE(en),
        .D(t290),
        .Q(t298),
        .R(reset)
    );
    (*LOC = "SLICE_X0Y6", BEL = "HFF"*)
    FDRE # (
        .INIT(1'b0),
        .IS_C_INVERTED(1'b0),
        .IS_D_INVERTED(1'b0),
        .IS_R_INVERTED(1'b0)
    ) __t299 (
        .C(clock),
        .CE(en),
        .D(t291),
        .Q(t299),
        .R(reset)
    );
    assign t89 = {t299, t298, t297, t296, t295, t294, t293, t292};
endmodule
