module main (
    input wire clock,
    input wire reset,
    input wire en,
    input wire [7:0] a0_0,
    input wire [7:0] a0_1,
    input wire [7:0] a0_2,
    input wire [7:0] a0_3,
    input wire [7:0] b0_0,
    input wire [7:0] b0_1,
    input wire [7:0] b0_2,
    input wire [7:0] b0_3,
    input wire [7:0] a1_0,
    input wire [7:0] a1_1,
    input wire [7:0] a1_2,
    input wire [7:0] a1_3,
    input wire [7:0] b1_0,
    input wire [7:0] b1_1,
    input wire [7:0] b1_2,
    input wire [7:0] b1_3,
    input wire [7:0] a2_0,
    input wire [7:0] a2_1,
    input wire [7:0] a2_2,
    input wire [7:0] a2_3,
    input wire [7:0] b2_0,
    input wire [7:0] b2_1,
    input wire [7:0] b2_2,
    input wire [7:0] b2_3,
    input wire [7:0] a3_0,
    input wire [7:0] a3_1,
    input wire [7:0] a3_2,
    input wire [7:0] a3_3,
    input wire [7:0] b3_0,
    input wire [7:0] b3_1,
    input wire [7:0] b3_2,
    input wire [7:0] b3_3,
    input wire [7:0] a4_0,
    input wire [7:0] a4_1,
    input wire [7:0] a4_2,
    input wire [7:0] a4_3,
    input wire [7:0] b4_0,
    input wire [7:0] b4_1,
    input wire [7:0] b4_2,
    input wire [7:0] b4_3,
    input wire [7:0] a5_0,
    input wire [7:0] a5_1,
    input wire [7:0] a5_2,
    input wire [7:0] a5_3,
    input wire [7:0] b5_0,
    input wire [7:0] b5_1,
    input wire [7:0] b5_2,
    input wire [7:0] b5_3,
    input wire [7:0] a6_0,
    input wire [7:0] a6_1,
    input wire [7:0] a6_2,
    input wire [7:0] a6_3,
    input wire [7:0] b6_0,
    input wire [7:0] b6_1,
    input wire [7:0] b6_2,
    input wire [7:0] b6_3,
    input wire [7:0] a7_0,
    input wire [7:0] a7_1,
    input wire [7:0] a7_2,
    input wire [7:0] a7_3,
    input wire [7:0] b7_0,
    input wire [7:0] b7_1,
    input wire [7:0] b7_2,
    input wire [7:0] b7_3,
    input wire [7:0] a8_0,
    input wire [7:0] a8_1,
    input wire [7:0] a8_2,
    input wire [7:0] a8_3,
    input wire [7:0] b8_0,
    input wire [7:0] b8_1,
    input wire [7:0] b8_2,
    input wire [7:0] b8_3,
    input wire [7:0] a9_0,
    input wire [7:0] a9_1,
    input wire [7:0] a9_2,
    input wire [7:0] a9_3,
    input wire [7:0] b9_0,
    input wire [7:0] b9_1,
    input wire [7:0] b9_2,
    input wire [7:0] b9_3,
    input wire [7:0] a10_0,
    input wire [7:0] a10_1,
    input wire [7:0] a10_2,
    input wire [7:0] a10_3,
    input wire [7:0] b10_0,
    input wire [7:0] b10_1,
    input wire [7:0] b10_2,
    input wire [7:0] b10_3,
    input wire [7:0] a11_0,
    input wire [7:0] a11_1,
    input wire [7:0] a11_2,
    input wire [7:0] a11_3,
    input wire [7:0] b11_0,
    input wire [7:0] b11_1,
    input wire [7:0] b11_2,
    input wire [7:0] b11_3,
    input wire [7:0] a12_0,
    input wire [7:0] a12_1,
    input wire [7:0] a12_2,
    input wire [7:0] a12_3,
    input wire [7:0] b12_0,
    input wire [7:0] b12_1,
    input wire [7:0] b12_2,
    input wire [7:0] b12_3,
    input wire [7:0] a13_0,
    input wire [7:0] a13_1,
    input wire [7:0] a13_2,
    input wire [7:0] a13_3,
    input wire [7:0] b13_0,
    input wire [7:0] b13_1,
    input wire [7:0] b13_2,
    input wire [7:0] b13_3,
    input wire [7:0] a14_0,
    input wire [7:0] a14_1,
    input wire [7:0] a14_2,
    input wire [7:0] a14_3,
    input wire [7:0] b14_0,
    input wire [7:0] b14_1,
    input wire [7:0] b14_2,
    input wire [7:0] b14_3,
    input wire [7:0] a15_0,
    input wire [7:0] a15_1,
    input wire [7:0] a15_2,
    input wire [7:0] a15_3,
    input wire [7:0] b15_0,
    input wire [7:0] b15_1,
    input wire [7:0] b15_2,
    input wire [7:0] b15_3,
    input wire [7:0] a16_0,
    input wire [7:0] a16_1,
    input wire [7:0] a16_2,
    input wire [7:0] a16_3,
    input wire [7:0] b16_0,
    input wire [7:0] b16_1,
    input wire [7:0] b16_2,
    input wire [7:0] b16_3,
    input wire [7:0] a17_0,
    input wire [7:0] a17_1,
    input wire [7:0] a17_2,
    input wire [7:0] a17_3,
    input wire [7:0] b17_0,
    input wire [7:0] b17_1,
    input wire [7:0] b17_2,
    input wire [7:0] b17_3,
    input wire [7:0] a18_0,
    input wire [7:0] a18_1,
    input wire [7:0] a18_2,
    input wire [7:0] a18_3,
    input wire [7:0] b18_0,
    input wire [7:0] b18_1,
    input wire [7:0] b18_2,
    input wire [7:0] b18_3,
    input wire [7:0] a19_0,
    input wire [7:0] a19_1,
    input wire [7:0] a19_2,
    input wire [7:0] a19_3,
    input wire [7:0] b19_0,
    input wire [7:0] b19_1,
    input wire [7:0] b19_2,
    input wire [7:0] b19_3,
    input wire [7:0] a20_0,
    input wire [7:0] a20_1,
    input wire [7:0] a20_2,
    input wire [7:0] a20_3,
    input wire [7:0] b20_0,
    input wire [7:0] b20_1,
    input wire [7:0] b20_2,
    input wire [7:0] b20_3,
    input wire [7:0] a21_0,
    input wire [7:0] a21_1,
    input wire [7:0] a21_2,
    input wire [7:0] a21_3,
    input wire [7:0] b21_0,
    input wire [7:0] b21_1,
    input wire [7:0] b21_2,
    input wire [7:0] b21_3,
    input wire [7:0] a22_0,
    input wire [7:0] a22_1,
    input wire [7:0] a22_2,
    input wire [7:0] a22_3,
    input wire [7:0] b22_0,
    input wire [7:0] b22_1,
    input wire [7:0] b22_2,
    input wire [7:0] b22_3,
    input wire [7:0] a23_0,
    input wire [7:0] a23_1,
    input wire [7:0] a23_2,
    input wire [7:0] a23_3,
    input wire [7:0] b23_0,
    input wire [7:0] b23_1,
    input wire [7:0] b23_2,
    input wire [7:0] b23_3,
    input wire [7:0] a24_0,
    input wire [7:0] a24_1,
    input wire [7:0] a24_2,
    input wire [7:0] a24_3,
    input wire [7:0] b24_0,
    input wire [7:0] b24_1,
    input wire [7:0] b24_2,
    input wire [7:0] b24_3,
    input wire [7:0] a25_0,
    input wire [7:0] a25_1,
    input wire [7:0] a25_2,
    input wire [7:0] a25_3,
    input wire [7:0] b25_0,
    input wire [7:0] b25_1,
    input wire [7:0] b25_2,
    input wire [7:0] b25_3,
    input wire [7:0] a26_0,
    input wire [7:0] a26_1,
    input wire [7:0] a26_2,
    input wire [7:0] a26_3,
    input wire [7:0] b26_0,
    input wire [7:0] b26_1,
    input wire [7:0] b26_2,
    input wire [7:0] b26_3,
    input wire [7:0] a27_0,
    input wire [7:0] a27_1,
    input wire [7:0] a27_2,
    input wire [7:0] a27_3,
    input wire [7:0] b27_0,
    input wire [7:0] b27_1,
    input wire [7:0] b27_2,
    input wire [7:0] b27_3,
    input wire [7:0] a28_0,
    input wire [7:0] a28_1,
    input wire [7:0] a28_2,
    input wire [7:0] a28_3,
    input wire [7:0] b28_0,
    input wire [7:0] b28_1,
    input wire [7:0] b28_2,
    input wire [7:0] b28_3,
    input wire [7:0] a29_0,
    input wire [7:0] a29_1,
    input wire [7:0] a29_2,
    input wire [7:0] a29_3,
    input wire [7:0] b29_0,
    input wire [7:0] b29_1,
    input wire [7:0] b29_2,
    input wire [7:0] b29_3,
    input wire [7:0] a30_0,
    input wire [7:0] a30_1,
    input wire [7:0] a30_2,
    input wire [7:0] a30_3,
    input wire [7:0] b30_0,
    input wire [7:0] b30_1,
    input wire [7:0] b30_2,
    input wire [7:0] b30_3,
    input wire [7:0] a31_0,
    input wire [7:0] a31_1,
    input wire [7:0] a31_2,
    input wire [7:0] a31_3,
    input wire [7:0] b31_0,
    input wire [7:0] b31_1,
    input wire [7:0] b31_2,
    input wire [7:0] b31_3,
    input wire [7:0] a32_0,
    input wire [7:0] a32_1,
    input wire [7:0] a32_2,
    input wire [7:0] a32_3,
    input wire [7:0] b32_0,
    input wire [7:0] b32_1,
    input wire [7:0] b32_2,
    input wire [7:0] b32_3,
    input wire [7:0] a33_0,
    input wire [7:0] a33_1,
    input wire [7:0] a33_2,
    input wire [7:0] a33_3,
    input wire [7:0] b33_0,
    input wire [7:0] b33_1,
    input wire [7:0] b33_2,
    input wire [7:0] b33_3,
    input wire [7:0] a34_0,
    input wire [7:0] a34_1,
    input wire [7:0] a34_2,
    input wire [7:0] a34_3,
    input wire [7:0] b34_0,
    input wire [7:0] b34_1,
    input wire [7:0] b34_2,
    input wire [7:0] b34_3,
    input wire [7:0] a35_0,
    input wire [7:0] a35_1,
    input wire [7:0] a35_2,
    input wire [7:0] a35_3,
    input wire [7:0] b35_0,
    input wire [7:0] b35_1,
    input wire [7:0] b35_2,
    input wire [7:0] b35_3,
    input wire [7:0] a36_0,
    input wire [7:0] a36_1,
    input wire [7:0] a36_2,
    input wire [7:0] a36_3,
    input wire [7:0] b36_0,
    input wire [7:0] b36_1,
    input wire [7:0] b36_2,
    input wire [7:0] b36_3,
    input wire [7:0] a37_0,
    input wire [7:0] a37_1,
    input wire [7:0] a37_2,
    input wire [7:0] a37_3,
    input wire [7:0] b37_0,
    input wire [7:0] b37_1,
    input wire [7:0] b37_2,
    input wire [7:0] b37_3,
    input wire [7:0] a38_0,
    input wire [7:0] a38_1,
    input wire [7:0] a38_2,
    input wire [7:0] a38_3,
    input wire [7:0] b38_0,
    input wire [7:0] b38_1,
    input wire [7:0] b38_2,
    input wire [7:0] b38_3,
    input wire [7:0] a39_0,
    input wire [7:0] a39_1,
    input wire [7:0] a39_2,
    input wire [7:0] a39_3,
    input wire [7:0] b39_0,
    input wire [7:0] b39_1,
    input wire [7:0] b39_2,
    input wire [7:0] b39_3,
    input wire [7:0] a40_0,
    input wire [7:0] a40_1,
    input wire [7:0] a40_2,
    input wire [7:0] a40_3,
    input wire [7:0] b40_0,
    input wire [7:0] b40_1,
    input wire [7:0] b40_2,
    input wire [7:0] b40_3,
    input wire [7:0] a41_0,
    input wire [7:0] a41_1,
    input wire [7:0] a41_2,
    input wire [7:0] a41_3,
    input wire [7:0] b41_0,
    input wire [7:0] b41_1,
    input wire [7:0] b41_2,
    input wire [7:0] b41_3,
    input wire [7:0] a42_0,
    input wire [7:0] a42_1,
    input wire [7:0] a42_2,
    input wire [7:0] a42_3,
    input wire [7:0] b42_0,
    input wire [7:0] b42_1,
    input wire [7:0] b42_2,
    input wire [7:0] b42_3,
    input wire [7:0] a43_0,
    input wire [7:0] a43_1,
    input wire [7:0] a43_2,
    input wire [7:0] a43_3,
    input wire [7:0] b43_0,
    input wire [7:0] b43_1,
    input wire [7:0] b43_2,
    input wire [7:0] b43_3,
    input wire [7:0] a44_0,
    input wire [7:0] a44_1,
    input wire [7:0] a44_2,
    input wire [7:0] a44_3,
    input wire [7:0] b44_0,
    input wire [7:0] b44_1,
    input wire [7:0] b44_2,
    input wire [7:0] b44_3,
    input wire [7:0] a45_0,
    input wire [7:0] a45_1,
    input wire [7:0] a45_2,
    input wire [7:0] a45_3,
    input wire [7:0] b45_0,
    input wire [7:0] b45_1,
    input wire [7:0] b45_2,
    input wire [7:0] b45_3,
    input wire [7:0] a46_0,
    input wire [7:0] a46_1,
    input wire [7:0] a46_2,
    input wire [7:0] a46_3,
    input wire [7:0] b46_0,
    input wire [7:0] b46_1,
    input wire [7:0] b46_2,
    input wire [7:0] b46_3,
    input wire [7:0] a47_0,
    input wire [7:0] a47_1,
    input wire [7:0] a47_2,
    input wire [7:0] a47_3,
    input wire [7:0] b47_0,
    input wire [7:0] b47_1,
    input wire [7:0] b47_2,
    input wire [7:0] b47_3,
    input wire [7:0] a48_0,
    input wire [7:0] a48_1,
    input wire [7:0] a48_2,
    input wire [7:0] a48_3,
    input wire [7:0] b48_0,
    input wire [7:0] b48_1,
    input wire [7:0] b48_2,
    input wire [7:0] b48_3,
    input wire [7:0] a49_0,
    input wire [7:0] a49_1,
    input wire [7:0] a49_2,
    input wire [7:0] a49_3,
    input wire [7:0] b49_0,
    input wire [7:0] b49_1,
    input wire [7:0] b49_2,
    input wire [7:0] b49_3,
    input wire [7:0] a50_0,
    input wire [7:0] a50_1,
    input wire [7:0] a50_2,
    input wire [7:0] a50_3,
    input wire [7:0] b50_0,
    input wire [7:0] b50_1,
    input wire [7:0] b50_2,
    input wire [7:0] b50_3,
    input wire [7:0] a51_0,
    input wire [7:0] a51_1,
    input wire [7:0] a51_2,
    input wire [7:0] a51_3,
    input wire [7:0] b51_0,
    input wire [7:0] b51_1,
    input wire [7:0] b51_2,
    input wire [7:0] b51_3,
    input wire [7:0] a52_0,
    input wire [7:0] a52_1,
    input wire [7:0] a52_2,
    input wire [7:0] a52_3,
    input wire [7:0] b52_0,
    input wire [7:0] b52_1,
    input wire [7:0] b52_2,
    input wire [7:0] b52_3,
    input wire [7:0] a53_0,
    input wire [7:0] a53_1,
    input wire [7:0] a53_2,
    input wire [7:0] a53_3,
    input wire [7:0] b53_0,
    input wire [7:0] b53_1,
    input wire [7:0] b53_2,
    input wire [7:0] b53_3,
    input wire [7:0] a54_0,
    input wire [7:0] a54_1,
    input wire [7:0] a54_2,
    input wire [7:0] a54_3,
    input wire [7:0] b54_0,
    input wire [7:0] b54_1,
    input wire [7:0] b54_2,
    input wire [7:0] b54_3,
    input wire [7:0] a55_0,
    input wire [7:0] a55_1,
    input wire [7:0] a55_2,
    input wire [7:0] a55_3,
    input wire [7:0] b55_0,
    input wire [7:0] b55_1,
    input wire [7:0] b55_2,
    input wire [7:0] b55_3,
    input wire [7:0] a56_0,
    input wire [7:0] a56_1,
    input wire [7:0] a56_2,
    input wire [7:0] a56_3,
    input wire [7:0] b56_0,
    input wire [7:0] b56_1,
    input wire [7:0] b56_2,
    input wire [7:0] b56_3,
    input wire [7:0] a57_0,
    input wire [7:0] a57_1,
    input wire [7:0] a57_2,
    input wire [7:0] a57_3,
    input wire [7:0] b57_0,
    input wire [7:0] b57_1,
    input wire [7:0] b57_2,
    input wire [7:0] b57_3,
    input wire [7:0] a58_0,
    input wire [7:0] a58_1,
    input wire [7:0] a58_2,
    input wire [7:0] a58_3,
    input wire [7:0] b58_0,
    input wire [7:0] b58_1,
    input wire [7:0] b58_2,
    input wire [7:0] b58_3,
    input wire [7:0] a59_0,
    input wire [7:0] a59_1,
    input wire [7:0] a59_2,
    input wire [7:0] a59_3,
    input wire [7:0] b59_0,
    input wire [7:0] b59_1,
    input wire [7:0] b59_2,
    input wire [7:0] b59_3,
    input wire [7:0] a60_0,
    input wire [7:0] a60_1,
    input wire [7:0] a60_2,
    input wire [7:0] a60_3,
    input wire [7:0] b60_0,
    input wire [7:0] b60_1,
    input wire [7:0] b60_2,
    input wire [7:0] b60_3,
    input wire [7:0] a61_0,
    input wire [7:0] a61_1,
    input wire [7:0] a61_2,
    input wire [7:0] a61_3,
    input wire [7:0] b61_0,
    input wire [7:0] b61_1,
    input wire [7:0] b61_2,
    input wire [7:0] b61_3,
    input wire [7:0] a62_0,
    input wire [7:0] a62_1,
    input wire [7:0] a62_2,
    input wire [7:0] a62_3,
    input wire [7:0] b62_0,
    input wire [7:0] b62_1,
    input wire [7:0] b62_2,
    input wire [7:0] b62_3,
    input wire [7:0] a63_0,
    input wire [7:0] a63_1,
    input wire [7:0] a63_2,
    input wire [7:0] a63_3,
    input wire [7:0] b63_0,
    input wire [7:0] b63_1,
    input wire [7:0] b63_2,
    input wire [7:0] b63_3,
    input wire [7:0] a64_0,
    input wire [7:0] a64_1,
    input wire [7:0] a64_2,
    input wire [7:0] a64_3,
    input wire [7:0] b64_0,
    input wire [7:0] b64_1,
    input wire [7:0] b64_2,
    input wire [7:0] b64_3,
    input wire [7:0] a65_0,
    input wire [7:0] a65_1,
    input wire [7:0] a65_2,
    input wire [7:0] a65_3,
    input wire [7:0] b65_0,
    input wire [7:0] b65_1,
    input wire [7:0] b65_2,
    input wire [7:0] b65_3,
    input wire [7:0] a66_0,
    input wire [7:0] a66_1,
    input wire [7:0] a66_2,
    input wire [7:0] a66_3,
    input wire [7:0] b66_0,
    input wire [7:0] b66_1,
    input wire [7:0] b66_2,
    input wire [7:0] b66_3,
    input wire [7:0] a67_0,
    input wire [7:0] a67_1,
    input wire [7:0] a67_2,
    input wire [7:0] a67_3,
    input wire [7:0] b67_0,
    input wire [7:0] b67_1,
    input wire [7:0] b67_2,
    input wire [7:0] b67_3,
    input wire [7:0] a68_0,
    input wire [7:0] a68_1,
    input wire [7:0] a68_2,
    input wire [7:0] a68_3,
    input wire [7:0] b68_0,
    input wire [7:0] b68_1,
    input wire [7:0] b68_2,
    input wire [7:0] b68_3,
    input wire [7:0] a69_0,
    input wire [7:0] a69_1,
    input wire [7:0] a69_2,
    input wire [7:0] a69_3,
    input wire [7:0] b69_0,
    input wire [7:0] b69_1,
    input wire [7:0] b69_2,
    input wire [7:0] b69_3,
    input wire [7:0] a70_0,
    input wire [7:0] a70_1,
    input wire [7:0] a70_2,
    input wire [7:0] a70_3,
    input wire [7:0] b70_0,
    input wire [7:0] b70_1,
    input wire [7:0] b70_2,
    input wire [7:0] b70_3,
    input wire [7:0] a71_0,
    input wire [7:0] a71_1,
    input wire [7:0] a71_2,
    input wire [7:0] a71_3,
    input wire [7:0] b71_0,
    input wire [7:0] b71_1,
    input wire [7:0] b71_2,
    input wire [7:0] b71_3,
    input wire [7:0] a72_0,
    input wire [7:0] a72_1,
    input wire [7:0] a72_2,
    input wire [7:0] a72_3,
    input wire [7:0] b72_0,
    input wire [7:0] b72_1,
    input wire [7:0] b72_2,
    input wire [7:0] b72_3,
    input wire [7:0] a73_0,
    input wire [7:0] a73_1,
    input wire [7:0] a73_2,
    input wire [7:0] a73_3,
    input wire [7:0] b73_0,
    input wire [7:0] b73_1,
    input wire [7:0] b73_2,
    input wire [7:0] b73_3,
    input wire [7:0] a74_0,
    input wire [7:0] a74_1,
    input wire [7:0] a74_2,
    input wire [7:0] a74_3,
    input wire [7:0] b74_0,
    input wire [7:0] b74_1,
    input wire [7:0] b74_2,
    input wire [7:0] b74_3,
    input wire [7:0] a75_0,
    input wire [7:0] a75_1,
    input wire [7:0] a75_2,
    input wire [7:0] a75_3,
    input wire [7:0] b75_0,
    input wire [7:0] b75_1,
    input wire [7:0] b75_2,
    input wire [7:0] b75_3,
    input wire [7:0] a76_0,
    input wire [7:0] a76_1,
    input wire [7:0] a76_2,
    input wire [7:0] a76_3,
    input wire [7:0] b76_0,
    input wire [7:0] b76_1,
    input wire [7:0] b76_2,
    input wire [7:0] b76_3,
    input wire [7:0] a77_0,
    input wire [7:0] a77_1,
    input wire [7:0] a77_2,
    input wire [7:0] a77_3,
    input wire [7:0] b77_0,
    input wire [7:0] b77_1,
    input wire [7:0] b77_2,
    input wire [7:0] b77_3,
    input wire [7:0] a78_0,
    input wire [7:0] a78_1,
    input wire [7:0] a78_2,
    input wire [7:0] a78_3,
    input wire [7:0] b78_0,
    input wire [7:0] b78_1,
    input wire [7:0] b78_2,
    input wire [7:0] b78_3,
    input wire [7:0] a79_0,
    input wire [7:0] a79_1,
    input wire [7:0] a79_2,
    input wire [7:0] a79_3,
    input wire [7:0] b79_0,
    input wire [7:0] b79_1,
    input wire [7:0] b79_2,
    input wire [7:0] b79_3,
    input wire [7:0] a80_0,
    input wire [7:0] a80_1,
    input wire [7:0] a80_2,
    input wire [7:0] a80_3,
    input wire [7:0] b80_0,
    input wire [7:0] b80_1,
    input wire [7:0] b80_2,
    input wire [7:0] b80_3,
    input wire [7:0] a81_0,
    input wire [7:0] a81_1,
    input wire [7:0] a81_2,
    input wire [7:0] a81_3,
    input wire [7:0] b81_0,
    input wire [7:0] b81_1,
    input wire [7:0] b81_2,
    input wire [7:0] b81_3,
    input wire [7:0] a82_0,
    input wire [7:0] a82_1,
    input wire [7:0] a82_2,
    input wire [7:0] a82_3,
    input wire [7:0] b82_0,
    input wire [7:0] b82_1,
    input wire [7:0] b82_2,
    input wire [7:0] b82_3,
    input wire [7:0] a83_0,
    input wire [7:0] a83_1,
    input wire [7:0] a83_2,
    input wire [7:0] a83_3,
    input wire [7:0] b83_0,
    input wire [7:0] b83_1,
    input wire [7:0] b83_2,
    input wire [7:0] b83_3,
    input wire [7:0] a84_0,
    input wire [7:0] a84_1,
    input wire [7:0] a84_2,
    input wire [7:0] a84_3,
    input wire [7:0] b84_0,
    input wire [7:0] b84_1,
    input wire [7:0] b84_2,
    input wire [7:0] b84_3,
    input wire [7:0] a85_0,
    input wire [7:0] a85_1,
    input wire [7:0] a85_2,
    input wire [7:0] a85_3,
    input wire [7:0] b85_0,
    input wire [7:0] b85_1,
    input wire [7:0] b85_2,
    input wire [7:0] b85_3,
    input wire [7:0] a86_0,
    input wire [7:0] a86_1,
    input wire [7:0] a86_2,
    input wire [7:0] a86_3,
    input wire [7:0] b86_0,
    input wire [7:0] b86_1,
    input wire [7:0] b86_2,
    input wire [7:0] b86_3,
    input wire [7:0] a87_0,
    input wire [7:0] a87_1,
    input wire [7:0] a87_2,
    input wire [7:0] a87_3,
    input wire [7:0] b87_0,
    input wire [7:0] b87_1,
    input wire [7:0] b87_2,
    input wire [7:0] b87_3,
    input wire [7:0] a88_0,
    input wire [7:0] a88_1,
    input wire [7:0] a88_2,
    input wire [7:0] a88_3,
    input wire [7:0] b88_0,
    input wire [7:0] b88_1,
    input wire [7:0] b88_2,
    input wire [7:0] b88_3,
    input wire [7:0] a89_0,
    input wire [7:0] a89_1,
    input wire [7:0] a89_2,
    input wire [7:0] a89_3,
    input wire [7:0] b89_0,
    input wire [7:0] b89_1,
    input wire [7:0] b89_2,
    input wire [7:0] b89_3,
    input wire [7:0] a90_0,
    input wire [7:0] a90_1,
    input wire [7:0] a90_2,
    input wire [7:0] a90_3,
    input wire [7:0] b90_0,
    input wire [7:0] b90_1,
    input wire [7:0] b90_2,
    input wire [7:0] b90_3,
    input wire [7:0] a91_0,
    input wire [7:0] a91_1,
    input wire [7:0] a91_2,
    input wire [7:0] a91_3,
    input wire [7:0] b91_0,
    input wire [7:0] b91_1,
    input wire [7:0] b91_2,
    input wire [7:0] b91_3,
    input wire [7:0] a92_0,
    input wire [7:0] a92_1,
    input wire [7:0] a92_2,
    input wire [7:0] a92_3,
    input wire [7:0] b92_0,
    input wire [7:0] b92_1,
    input wire [7:0] b92_2,
    input wire [7:0] b92_3,
    input wire [7:0] a93_0,
    input wire [7:0] a93_1,
    input wire [7:0] a93_2,
    input wire [7:0] a93_3,
    input wire [7:0] b93_0,
    input wire [7:0] b93_1,
    input wire [7:0] b93_2,
    input wire [7:0] b93_3,
    input wire [7:0] a94_0,
    input wire [7:0] a94_1,
    input wire [7:0] a94_2,
    input wire [7:0] a94_3,
    input wire [7:0] b94_0,
    input wire [7:0] b94_1,
    input wire [7:0] b94_2,
    input wire [7:0] b94_3,
    input wire [7:0] a95_0,
    input wire [7:0] a95_1,
    input wire [7:0] a95_2,
    input wire [7:0] a95_3,
    input wire [7:0] b95_0,
    input wire [7:0] b95_1,
    input wire [7:0] b95_2,
    input wire [7:0] b95_3,
    input wire [7:0] a96_0,
    input wire [7:0] a96_1,
    input wire [7:0] a96_2,
    input wire [7:0] a96_3,
    input wire [7:0] b96_0,
    input wire [7:0] b96_1,
    input wire [7:0] b96_2,
    input wire [7:0] b96_3,
    input wire [7:0] a97_0,
    input wire [7:0] a97_1,
    input wire [7:0] a97_2,
    input wire [7:0] a97_3,
    input wire [7:0] b97_0,
    input wire [7:0] b97_1,
    input wire [7:0] b97_2,
    input wire [7:0] b97_3,
    input wire [7:0] a98_0,
    input wire [7:0] a98_1,
    input wire [7:0] a98_2,
    input wire [7:0] a98_3,
    input wire [7:0] b98_0,
    input wire [7:0] b98_1,
    input wire [7:0] b98_2,
    input wire [7:0] b98_3,
    input wire [7:0] a99_0,
    input wire [7:0] a99_1,
    input wire [7:0] a99_2,
    input wire [7:0] a99_3,
    input wire [7:0] b99_0,
    input wire [7:0] b99_1,
    input wire [7:0] b99_2,
    input wire [7:0] b99_3,
    input wire [7:0] a100_0,
    input wire [7:0] a100_1,
    input wire [7:0] a100_2,
    input wire [7:0] a100_3,
    input wire [7:0] b100_0,
    input wire [7:0] b100_1,
    input wire [7:0] b100_2,
    input wire [7:0] b100_3,
    input wire [7:0] a101_0,
    input wire [7:0] a101_1,
    input wire [7:0] a101_2,
    input wire [7:0] a101_3,
    input wire [7:0] b101_0,
    input wire [7:0] b101_1,
    input wire [7:0] b101_2,
    input wire [7:0] b101_3,
    input wire [7:0] a102_0,
    input wire [7:0] a102_1,
    input wire [7:0] a102_2,
    input wire [7:0] a102_3,
    input wire [7:0] b102_0,
    input wire [7:0] b102_1,
    input wire [7:0] b102_2,
    input wire [7:0] b102_3,
    input wire [7:0] a103_0,
    input wire [7:0] a103_1,
    input wire [7:0] a103_2,
    input wire [7:0] a103_3,
    input wire [7:0] b103_0,
    input wire [7:0] b103_1,
    input wire [7:0] b103_2,
    input wire [7:0] b103_3,
    input wire [7:0] a104_0,
    input wire [7:0] a104_1,
    input wire [7:0] a104_2,
    input wire [7:0] a104_3,
    input wire [7:0] b104_0,
    input wire [7:0] b104_1,
    input wire [7:0] b104_2,
    input wire [7:0] b104_3,
    input wire [7:0] a105_0,
    input wire [7:0] a105_1,
    input wire [7:0] a105_2,
    input wire [7:0] a105_3,
    input wire [7:0] b105_0,
    input wire [7:0] b105_1,
    input wire [7:0] b105_2,
    input wire [7:0] b105_3,
    input wire [7:0] a106_0,
    input wire [7:0] a106_1,
    input wire [7:0] a106_2,
    input wire [7:0] a106_3,
    input wire [7:0] b106_0,
    input wire [7:0] b106_1,
    input wire [7:0] b106_2,
    input wire [7:0] b106_3,
    input wire [7:0] a107_0,
    input wire [7:0] a107_1,
    input wire [7:0] a107_2,
    input wire [7:0] a107_3,
    input wire [7:0] b107_0,
    input wire [7:0] b107_1,
    input wire [7:0] b107_2,
    input wire [7:0] b107_3,
    input wire [7:0] a108_0,
    input wire [7:0] a108_1,
    input wire [7:0] a108_2,
    input wire [7:0] a108_3,
    input wire [7:0] b108_0,
    input wire [7:0] b108_1,
    input wire [7:0] b108_2,
    input wire [7:0] b108_3,
    input wire [7:0] a109_0,
    input wire [7:0] a109_1,
    input wire [7:0] a109_2,
    input wire [7:0] a109_3,
    input wire [7:0] b109_0,
    input wire [7:0] b109_1,
    input wire [7:0] b109_2,
    input wire [7:0] b109_3,
    input wire [7:0] a110_0,
    input wire [7:0] a110_1,
    input wire [7:0] a110_2,
    input wire [7:0] a110_3,
    input wire [7:0] b110_0,
    input wire [7:0] b110_1,
    input wire [7:0] b110_2,
    input wire [7:0] b110_3,
    input wire [7:0] a111_0,
    input wire [7:0] a111_1,
    input wire [7:0] a111_2,
    input wire [7:0] a111_3,
    input wire [7:0] b111_0,
    input wire [7:0] b111_1,
    input wire [7:0] b111_2,
    input wire [7:0] b111_3,
    input wire [7:0] a112_0,
    input wire [7:0] a112_1,
    input wire [7:0] a112_2,
    input wire [7:0] a112_3,
    input wire [7:0] b112_0,
    input wire [7:0] b112_1,
    input wire [7:0] b112_2,
    input wire [7:0] b112_3,
    input wire [7:0] a113_0,
    input wire [7:0] a113_1,
    input wire [7:0] a113_2,
    input wire [7:0] a113_3,
    input wire [7:0] b113_0,
    input wire [7:0] b113_1,
    input wire [7:0] b113_2,
    input wire [7:0] b113_3,
    input wire [7:0] a114_0,
    input wire [7:0] a114_1,
    input wire [7:0] a114_2,
    input wire [7:0] a114_3,
    input wire [7:0] b114_0,
    input wire [7:0] b114_1,
    input wire [7:0] b114_2,
    input wire [7:0] b114_3,
    input wire [7:0] a115_0,
    input wire [7:0] a115_1,
    input wire [7:0] a115_2,
    input wire [7:0] a115_3,
    input wire [7:0] b115_0,
    input wire [7:0] b115_1,
    input wire [7:0] b115_2,
    input wire [7:0] b115_3,
    input wire [7:0] a116_0,
    input wire [7:0] a116_1,
    input wire [7:0] a116_2,
    input wire [7:0] a116_3,
    input wire [7:0] b116_0,
    input wire [7:0] b116_1,
    input wire [7:0] b116_2,
    input wire [7:0] b116_3,
    input wire [7:0] a117_0,
    input wire [7:0] a117_1,
    input wire [7:0] a117_2,
    input wire [7:0] a117_3,
    input wire [7:0] b117_0,
    input wire [7:0] b117_1,
    input wire [7:0] b117_2,
    input wire [7:0] b117_3,
    input wire [7:0] a118_0,
    input wire [7:0] a118_1,
    input wire [7:0] a118_2,
    input wire [7:0] a118_3,
    input wire [7:0] b118_0,
    input wire [7:0] b118_1,
    input wire [7:0] b118_2,
    input wire [7:0] b118_3,
    input wire [7:0] a119_0,
    input wire [7:0] a119_1,
    input wire [7:0] a119_2,
    input wire [7:0] a119_3,
    input wire [7:0] b119_0,
    input wire [7:0] b119_1,
    input wire [7:0] b119_2,
    input wire [7:0] b119_3,
    input wire [7:0] a120_0,
    input wire [7:0] a120_1,
    input wire [7:0] a120_2,
    input wire [7:0] a120_3,
    input wire [7:0] b120_0,
    input wire [7:0] b120_1,
    input wire [7:0] b120_2,
    input wire [7:0] b120_3,
    input wire [7:0] a121_0,
    input wire [7:0] a121_1,
    input wire [7:0] a121_2,
    input wire [7:0] a121_3,
    input wire [7:0] b121_0,
    input wire [7:0] b121_1,
    input wire [7:0] b121_2,
    input wire [7:0] b121_3,
    input wire [7:0] a122_0,
    input wire [7:0] a122_1,
    input wire [7:0] a122_2,
    input wire [7:0] a122_3,
    input wire [7:0] b122_0,
    input wire [7:0] b122_1,
    input wire [7:0] b122_2,
    input wire [7:0] b122_3,
    input wire [7:0] a123_0,
    input wire [7:0] a123_1,
    input wire [7:0] a123_2,
    input wire [7:0] a123_3,
    input wire [7:0] b123_0,
    input wire [7:0] b123_1,
    input wire [7:0] b123_2,
    input wire [7:0] b123_3,
    input wire [7:0] a124_0,
    input wire [7:0] a124_1,
    input wire [7:0] a124_2,
    input wire [7:0] a124_3,
    input wire [7:0] b124_0,
    input wire [7:0] b124_1,
    input wire [7:0] b124_2,
    input wire [7:0] b124_3,
    input wire [7:0] a125_0,
    input wire [7:0] a125_1,
    input wire [7:0] a125_2,
    input wire [7:0] a125_3,
    input wire [7:0] b125_0,
    input wire [7:0] b125_1,
    input wire [7:0] b125_2,
    input wire [7:0] b125_3,
    input wire [7:0] a126_0,
    input wire [7:0] a126_1,
    input wire [7:0] a126_2,
    input wire [7:0] a126_3,
    input wire [7:0] b126_0,
    input wire [7:0] b126_1,
    input wire [7:0] b126_2,
    input wire [7:0] b126_3,
    input wire [7:0] a127_0,
    input wire [7:0] a127_1,
    input wire [7:0] a127_2,
    input wire [7:0] a127_3,
    input wire [7:0] b127_0,
    input wire [7:0] b127_1,
    input wire [7:0] b127_2,
    input wire [7:0] b127_3,
    output wire [7:0] y0_0,
    output wire [7:0] y0_1,
    output wire [7:0] y0_2,
    output wire [7:0] y0_3,
    output wire [7:0] y1_0,
    output wire [7:0] y1_1,
    output wire [7:0] y1_2,
    output wire [7:0] y1_3,
    output wire [7:0] y2_0,
    output wire [7:0] y2_1,
    output wire [7:0] y2_2,
    output wire [7:0] y2_3,
    output wire [7:0] y3_0,
    output wire [7:0] y3_1,
    output wire [7:0] y3_2,
    output wire [7:0] y3_3,
    output wire [7:0] y4_0,
    output wire [7:0] y4_1,
    output wire [7:0] y4_2,
    output wire [7:0] y4_3,
    output wire [7:0] y5_0,
    output wire [7:0] y5_1,
    output wire [7:0] y5_2,
    output wire [7:0] y5_3,
    output wire [7:0] y6_0,
    output wire [7:0] y6_1,
    output wire [7:0] y6_2,
    output wire [7:0] y6_3,
    output wire [7:0] y7_0,
    output wire [7:0] y7_1,
    output wire [7:0] y7_2,
    output wire [7:0] y7_3,
    output wire [7:0] y8_0,
    output wire [7:0] y8_1,
    output wire [7:0] y8_2,
    output wire [7:0] y8_3,
    output wire [7:0] y9_0,
    output wire [7:0] y9_1,
    output wire [7:0] y9_2,
    output wire [7:0] y9_3,
    output wire [7:0] y10_0,
    output wire [7:0] y10_1,
    output wire [7:0] y10_2,
    output wire [7:0] y10_3,
    output wire [7:0] y11_0,
    output wire [7:0] y11_1,
    output wire [7:0] y11_2,
    output wire [7:0] y11_3,
    output wire [7:0] y12_0,
    output wire [7:0] y12_1,
    output wire [7:0] y12_2,
    output wire [7:0] y12_3,
    output wire [7:0] y13_0,
    output wire [7:0] y13_1,
    output wire [7:0] y13_2,
    output wire [7:0] y13_3,
    output wire [7:0] y14_0,
    output wire [7:0] y14_1,
    output wire [7:0] y14_2,
    output wire [7:0] y14_3,
    output wire [7:0] y15_0,
    output wire [7:0] y15_1,
    output wire [7:0] y15_2,
    output wire [7:0] y15_3,
    output wire [7:0] y16_0,
    output wire [7:0] y16_1,
    output wire [7:0] y16_2,
    output wire [7:0] y16_3,
    output wire [7:0] y17_0,
    output wire [7:0] y17_1,
    output wire [7:0] y17_2,
    output wire [7:0] y17_3,
    output wire [7:0] y18_0,
    output wire [7:0] y18_1,
    output wire [7:0] y18_2,
    output wire [7:0] y18_3,
    output wire [7:0] y19_0,
    output wire [7:0] y19_1,
    output wire [7:0] y19_2,
    output wire [7:0] y19_3,
    output wire [7:0] y20_0,
    output wire [7:0] y20_1,
    output wire [7:0] y20_2,
    output wire [7:0] y20_3,
    output wire [7:0] y21_0,
    output wire [7:0] y21_1,
    output wire [7:0] y21_2,
    output wire [7:0] y21_3,
    output wire [7:0] y22_0,
    output wire [7:0] y22_1,
    output wire [7:0] y22_2,
    output wire [7:0] y22_3,
    output wire [7:0] y23_0,
    output wire [7:0] y23_1,
    output wire [7:0] y23_2,
    output wire [7:0] y23_3,
    output wire [7:0] y24_0,
    output wire [7:0] y24_1,
    output wire [7:0] y24_2,
    output wire [7:0] y24_3,
    output wire [7:0] y25_0,
    output wire [7:0] y25_1,
    output wire [7:0] y25_2,
    output wire [7:0] y25_3,
    output wire [7:0] y26_0,
    output wire [7:0] y26_1,
    output wire [7:0] y26_2,
    output wire [7:0] y26_3,
    output wire [7:0] y27_0,
    output wire [7:0] y27_1,
    output wire [7:0] y27_2,
    output wire [7:0] y27_3,
    output wire [7:0] y28_0,
    output wire [7:0] y28_1,
    output wire [7:0] y28_2,
    output wire [7:0] y28_3,
    output wire [7:0] y29_0,
    output wire [7:0] y29_1,
    output wire [7:0] y29_2,
    output wire [7:0] y29_3,
    output wire [7:0] y30_0,
    output wire [7:0] y30_1,
    output wire [7:0] y30_2,
    output wire [7:0] y30_3,
    output wire [7:0] y31_0,
    output wire [7:0] y31_1,
    output wire [7:0] y31_2,
    output wire [7:0] y31_3,
    output wire [7:0] y32_0,
    output wire [7:0] y32_1,
    output wire [7:0] y32_2,
    output wire [7:0] y32_3,
    output wire [7:0] y33_0,
    output wire [7:0] y33_1,
    output wire [7:0] y33_2,
    output wire [7:0] y33_3,
    output wire [7:0] y34_0,
    output wire [7:0] y34_1,
    output wire [7:0] y34_2,
    output wire [7:0] y34_3,
    output wire [7:0] y35_0,
    output wire [7:0] y35_1,
    output wire [7:0] y35_2,
    output wire [7:0] y35_3,
    output wire [7:0] y36_0,
    output wire [7:0] y36_1,
    output wire [7:0] y36_2,
    output wire [7:0] y36_3,
    output wire [7:0] y37_0,
    output wire [7:0] y37_1,
    output wire [7:0] y37_2,
    output wire [7:0] y37_3,
    output wire [7:0] y38_0,
    output wire [7:0] y38_1,
    output wire [7:0] y38_2,
    output wire [7:0] y38_3,
    output wire [7:0] y39_0,
    output wire [7:0] y39_1,
    output wire [7:0] y39_2,
    output wire [7:0] y39_3,
    output wire [7:0] y40_0,
    output wire [7:0] y40_1,
    output wire [7:0] y40_2,
    output wire [7:0] y40_3,
    output wire [7:0] y41_0,
    output wire [7:0] y41_1,
    output wire [7:0] y41_2,
    output wire [7:0] y41_3,
    output wire [7:0] y42_0,
    output wire [7:0] y42_1,
    output wire [7:0] y42_2,
    output wire [7:0] y42_3,
    output wire [7:0] y43_0,
    output wire [7:0] y43_1,
    output wire [7:0] y43_2,
    output wire [7:0] y43_3,
    output wire [7:0] y44_0,
    output wire [7:0] y44_1,
    output wire [7:0] y44_2,
    output wire [7:0] y44_3,
    output wire [7:0] y45_0,
    output wire [7:0] y45_1,
    output wire [7:0] y45_2,
    output wire [7:0] y45_3,
    output wire [7:0] y46_0,
    output wire [7:0] y46_1,
    output wire [7:0] y46_2,
    output wire [7:0] y46_3,
    output wire [7:0] y47_0,
    output wire [7:0] y47_1,
    output wire [7:0] y47_2,
    output wire [7:0] y47_3,
    output wire [7:0] y48_0,
    output wire [7:0] y48_1,
    output wire [7:0] y48_2,
    output wire [7:0] y48_3,
    output wire [7:0] y49_0,
    output wire [7:0] y49_1,
    output wire [7:0] y49_2,
    output wire [7:0] y49_3,
    output wire [7:0] y50_0,
    output wire [7:0] y50_1,
    output wire [7:0] y50_2,
    output wire [7:0] y50_3,
    output wire [7:0] y51_0,
    output wire [7:0] y51_1,
    output wire [7:0] y51_2,
    output wire [7:0] y51_3,
    output wire [7:0] y52_0,
    output wire [7:0] y52_1,
    output wire [7:0] y52_2,
    output wire [7:0] y52_3,
    output wire [7:0] y53_0,
    output wire [7:0] y53_1,
    output wire [7:0] y53_2,
    output wire [7:0] y53_3,
    output wire [7:0] y54_0,
    output wire [7:0] y54_1,
    output wire [7:0] y54_2,
    output wire [7:0] y54_3,
    output wire [7:0] y55_0,
    output wire [7:0] y55_1,
    output wire [7:0] y55_2,
    output wire [7:0] y55_3,
    output wire [7:0] y56_0,
    output wire [7:0] y56_1,
    output wire [7:0] y56_2,
    output wire [7:0] y56_3,
    output wire [7:0] y57_0,
    output wire [7:0] y57_1,
    output wire [7:0] y57_2,
    output wire [7:0] y57_3,
    output wire [7:0] y58_0,
    output wire [7:0] y58_1,
    output wire [7:0] y58_2,
    output wire [7:0] y58_3,
    output wire [7:0] y59_0,
    output wire [7:0] y59_1,
    output wire [7:0] y59_2,
    output wire [7:0] y59_3,
    output wire [7:0] y60_0,
    output wire [7:0] y60_1,
    output wire [7:0] y60_2,
    output wire [7:0] y60_3,
    output wire [7:0] y61_0,
    output wire [7:0] y61_1,
    output wire [7:0] y61_2,
    output wire [7:0] y61_3,
    output wire [7:0] y62_0,
    output wire [7:0] y62_1,
    output wire [7:0] y62_2,
    output wire [7:0] y62_3,
    output wire [7:0] y63_0,
    output wire [7:0] y63_1,
    output wire [7:0] y63_2,
    output wire [7:0] y63_3,
    output wire [7:0] y64_0,
    output wire [7:0] y64_1,
    output wire [7:0] y64_2,
    output wire [7:0] y64_3,
    output wire [7:0] y65_0,
    output wire [7:0] y65_1,
    output wire [7:0] y65_2,
    output wire [7:0] y65_3,
    output wire [7:0] y66_0,
    output wire [7:0] y66_1,
    output wire [7:0] y66_2,
    output wire [7:0] y66_3,
    output wire [7:0] y67_0,
    output wire [7:0] y67_1,
    output wire [7:0] y67_2,
    output wire [7:0] y67_3,
    output wire [7:0] y68_0,
    output wire [7:0] y68_1,
    output wire [7:0] y68_2,
    output wire [7:0] y68_3,
    output wire [7:0] y69_0,
    output wire [7:0] y69_1,
    output wire [7:0] y69_2,
    output wire [7:0] y69_3,
    output wire [7:0] y70_0,
    output wire [7:0] y70_1,
    output wire [7:0] y70_2,
    output wire [7:0] y70_3,
    output wire [7:0] y71_0,
    output wire [7:0] y71_1,
    output wire [7:0] y71_2,
    output wire [7:0] y71_3,
    output wire [7:0] y72_0,
    output wire [7:0] y72_1,
    output wire [7:0] y72_2,
    output wire [7:0] y72_3,
    output wire [7:0] y73_0,
    output wire [7:0] y73_1,
    output wire [7:0] y73_2,
    output wire [7:0] y73_3,
    output wire [7:0] y74_0,
    output wire [7:0] y74_1,
    output wire [7:0] y74_2,
    output wire [7:0] y74_3,
    output wire [7:0] y75_0,
    output wire [7:0] y75_1,
    output wire [7:0] y75_2,
    output wire [7:0] y75_3,
    output wire [7:0] y76_0,
    output wire [7:0] y76_1,
    output wire [7:0] y76_2,
    output wire [7:0] y76_3,
    output wire [7:0] y77_0,
    output wire [7:0] y77_1,
    output wire [7:0] y77_2,
    output wire [7:0] y77_3,
    output wire [7:0] y78_0,
    output wire [7:0] y78_1,
    output wire [7:0] y78_2,
    output wire [7:0] y78_3,
    output wire [7:0] y79_0,
    output wire [7:0] y79_1,
    output wire [7:0] y79_2,
    output wire [7:0] y79_3,
    output wire [7:0] y80_0,
    output wire [7:0] y80_1,
    output wire [7:0] y80_2,
    output wire [7:0] y80_3,
    output wire [7:0] y81_0,
    output wire [7:0] y81_1,
    output wire [7:0] y81_2,
    output wire [7:0] y81_3,
    output wire [7:0] y82_0,
    output wire [7:0] y82_1,
    output wire [7:0] y82_2,
    output wire [7:0] y82_3,
    output wire [7:0] y83_0,
    output wire [7:0] y83_1,
    output wire [7:0] y83_2,
    output wire [7:0] y83_3,
    output wire [7:0] y84_0,
    output wire [7:0] y84_1,
    output wire [7:0] y84_2,
    output wire [7:0] y84_3,
    output wire [7:0] y85_0,
    output wire [7:0] y85_1,
    output wire [7:0] y85_2,
    output wire [7:0] y85_3,
    output wire [7:0] y86_0,
    output wire [7:0] y86_1,
    output wire [7:0] y86_2,
    output wire [7:0] y86_3,
    output wire [7:0] y87_0,
    output wire [7:0] y87_1,
    output wire [7:0] y87_2,
    output wire [7:0] y87_3,
    output wire [7:0] y88_0,
    output wire [7:0] y88_1,
    output wire [7:0] y88_2,
    output wire [7:0] y88_3,
    output wire [7:0] y89_0,
    output wire [7:0] y89_1,
    output wire [7:0] y89_2,
    output wire [7:0] y89_3,
    output wire [7:0] y90_0,
    output wire [7:0] y90_1,
    output wire [7:0] y90_2,
    output wire [7:0] y90_3,
    output wire [7:0] y91_0,
    output wire [7:0] y91_1,
    output wire [7:0] y91_2,
    output wire [7:0] y91_3,
    output wire [7:0] y92_0,
    output wire [7:0] y92_1,
    output wire [7:0] y92_2,
    output wire [7:0] y92_3,
    output wire [7:0] y93_0,
    output wire [7:0] y93_1,
    output wire [7:0] y93_2,
    output wire [7:0] y93_3,
    output wire [7:0] y94_0,
    output wire [7:0] y94_1,
    output wire [7:0] y94_2,
    output wire [7:0] y94_3,
    output wire [7:0] y95_0,
    output wire [7:0] y95_1,
    output wire [7:0] y95_2,
    output wire [7:0] y95_3,
    output wire [7:0] y96_0,
    output wire [7:0] y96_1,
    output wire [7:0] y96_2,
    output wire [7:0] y96_3,
    output wire [7:0] y97_0,
    output wire [7:0] y97_1,
    output wire [7:0] y97_2,
    output wire [7:0] y97_3,
    output wire [7:0] y98_0,
    output wire [7:0] y98_1,
    output wire [7:0] y98_2,
    output wire [7:0] y98_3,
    output wire [7:0] y99_0,
    output wire [7:0] y99_1,
    output wire [7:0] y99_2,
    output wire [7:0] y99_3,
    output wire [7:0] y100_0,
    output wire [7:0] y100_1,
    output wire [7:0] y100_2,
    output wire [7:0] y100_3,
    output wire [7:0] y101_0,
    output wire [7:0] y101_1,
    output wire [7:0] y101_2,
    output wire [7:0] y101_3,
    output wire [7:0] y102_0,
    output wire [7:0] y102_1,
    output wire [7:0] y102_2,
    output wire [7:0] y102_3,
    output wire [7:0] y103_0,
    output wire [7:0] y103_1,
    output wire [7:0] y103_2,
    output wire [7:0] y103_3,
    output wire [7:0] y104_0,
    output wire [7:0] y104_1,
    output wire [7:0] y104_2,
    output wire [7:0] y104_3,
    output wire [7:0] y105_0,
    output wire [7:0] y105_1,
    output wire [7:0] y105_2,
    output wire [7:0] y105_3,
    output wire [7:0] y106_0,
    output wire [7:0] y106_1,
    output wire [7:0] y106_2,
    output wire [7:0] y106_3,
    output wire [7:0] y107_0,
    output wire [7:0] y107_1,
    output wire [7:0] y107_2,
    output wire [7:0] y107_3,
    output wire [7:0] y108_0,
    output wire [7:0] y108_1,
    output wire [7:0] y108_2,
    output wire [7:0] y108_3,
    output wire [7:0] y109_0,
    output wire [7:0] y109_1,
    output wire [7:0] y109_2,
    output wire [7:0] y109_3,
    output wire [7:0] y110_0,
    output wire [7:0] y110_1,
    output wire [7:0] y110_2,
    output wire [7:0] y110_3,
    output wire [7:0] y111_0,
    output wire [7:0] y111_1,
    output wire [7:0] y111_2,
    output wire [7:0] y111_3,
    output wire [7:0] y112_0,
    output wire [7:0] y112_1,
    output wire [7:0] y112_2,
    output wire [7:0] y112_3,
    output wire [7:0] y113_0,
    output wire [7:0] y113_1,
    output wire [7:0] y113_2,
    output wire [7:0] y113_3,
    output wire [7:0] y114_0,
    output wire [7:0] y114_1,
    output wire [7:0] y114_2,
    output wire [7:0] y114_3,
    output wire [7:0] y115_0,
    output wire [7:0] y115_1,
    output wire [7:0] y115_2,
    output wire [7:0] y115_3,
    output wire [7:0] y116_0,
    output wire [7:0] y116_1,
    output wire [7:0] y116_2,
    output wire [7:0] y116_3,
    output wire [7:0] y117_0,
    output wire [7:0] y117_1,
    output wire [7:0] y117_2,
    output wire [7:0] y117_3,
    output wire [7:0] y118_0,
    output wire [7:0] y118_1,
    output wire [7:0] y118_2,
    output wire [7:0] y118_3,
    output wire [7:0] y119_0,
    output wire [7:0] y119_1,
    output wire [7:0] y119_2,
    output wire [7:0] y119_3,
    output wire [7:0] y120_0,
    output wire [7:0] y120_1,
    output wire [7:0] y120_2,
    output wire [7:0] y120_3,
    output wire [7:0] y121_0,
    output wire [7:0] y121_1,
    output wire [7:0] y121_2,
    output wire [7:0] y121_3,
    output wire [7:0] y122_0,
    output wire [7:0] y122_1,
    output wire [7:0] y122_2,
    output wire [7:0] y122_3,
    output wire [7:0] y123_0,
    output wire [7:0] y123_1,
    output wire [7:0] y123_2,
    output wire [7:0] y123_3,
    output wire [7:0] y124_0,
    output wire [7:0] y124_1,
    output wire [7:0] y124_2,
    output wire [7:0] y124_3,
    output wire [7:0] y125_0,
    output wire [7:0] y125_1,
    output wire [7:0] y125_2,
    output wire [7:0] y125_3,
    output wire [7:0] y126_0,
    output wire [7:0] y126_1,
    output wire [7:0] y126_2,
    output wire [7:0] y126_3,
    output wire [7:0] y127_0,
    output wire [7:0] y127_1,
    output wire [7:0] y127_2,
    output wire [7:0] y127_3
);
    wire gnd;
    wire vcc;
    wire [47:0] _y0;
    wire [47:0] _y1;
    wire [47:0] _y2;
    wire [47:0] _y3;
    wire [47:0] _y4;
    wire [47:0] _y5;
    wire [47:0] _y6;
    wire [47:0] _y7;
    wire [47:0] _y8;
    wire [47:0] _y9;
    wire [47:0] _y10;
    wire [47:0] _y11;
    wire [47:0] _y12;
    wire [47:0] _y13;
    wire [47:0] _y14;
    wire [47:0] _y15;
    wire [47:0] _y16;
    wire [47:0] _y17;
    wire [47:0] _y18;
    wire [47:0] _y19;
    wire [47:0] _y20;
    wire [47:0] _y21;
    wire [47:0] _y22;
    wire [47:0] _y23;
    wire [47:0] _y24;
    wire [47:0] _y25;
    wire [47:0] _y26;
    wire [47:0] _y27;
    wire [47:0] _y28;
    wire [47:0] _y29;
    wire [47:0] _y30;
    wire [47:0] _y31;
    wire [47:0] _y32;
    wire [47:0] _y33;
    wire [47:0] _y34;
    wire [47:0] _y35;
    wire [47:0] _y36;
    wire [47:0] _y37;
    wire [47:0] _y38;
    wire [47:0] _y39;
    wire [47:0] _y40;
    wire [47:0] _y41;
    wire [47:0] _y42;
    wire [47:0] _y43;
    wire [47:0] _y44;
    wire [47:0] _y45;
    wire [47:0] _y46;
    wire [47:0] _y47;
    wire [47:0] _y48;
    wire [47:0] _y49;
    wire [47:0] _y50;
    wire [47:0] _y51;
    wire [47:0] _y52;
    wire [47:0] _y53;
    wire [47:0] _y54;
    wire [47:0] _y55;
    wire [47:0] _y56;
    wire [47:0] _y57;
    wire [47:0] _y58;
    wire [47:0] _y59;
    wire [47:0] _y60;
    wire [47:0] _y61;
    wire [47:0] _y62;
    wire [47:0] _y63;
    wire [47:0] _y64;
    wire [47:0] _y65;
    wire [47:0] _y66;
    wire [47:0] _y67;
    wire [47:0] _y68;
    wire [47:0] _y69;
    wire [47:0] _y70;
    wire [47:0] _y71;
    wire [47:0] _y72;
    wire [47:0] _y73;
    wire [47:0] _y74;
    wire [47:0] _y75;
    wire [47:0] _y76;
    wire [47:0] _y77;
    wire [47:0] _y78;
    wire [47:0] _y79;
    wire [47:0] _y80;
    wire [47:0] _y81;
    wire [47:0] _y82;
    wire [47:0] _y83;
    wire [47:0] _y84;
    wire [47:0] _y85;
    wire [47:0] _y86;
    wire [47:0] _y87;
    wire [47:0] _y88;
    wire [47:0] _y89;
    wire [47:0] _y90;
    wire [47:0] _y91;
    wire [47:0] _y92;
    wire [47:0] _y93;
    wire [47:0] _y94;
    wire [47:0] _y95;
    wire [47:0] _y96;
    wire [47:0] _y97;
    wire [47:0] _y98;
    wire [47:0] _y99;
    wire [47:0] _y100;
    wire [47:0] _y101;
    wire [47:0] _y102;
    wire [47:0] _y103;
    wire [47:0] _y104;
    wire [47:0] _y105;
    wire [47:0] _y106;
    wire [47:0] _y107;
    wire [47:0] _y108;
    wire [47:0] _y109;
    wire [47:0] _y110;
    wire [47:0] _y111;
    wire [47:0] _y112;
    wire [47:0] _y113;
    wire [47:0] _y114;
    wire [47:0] _y115;
    wire [47:0] _y116;
    wire [47:0] _y117;
    wire [47:0] _y118;
    wire [47:0] _y119;
    wire [47:0] _y120;
    wire [47:0] _y121;
    wire [47:0] _y122;
    wire [47:0] _y123;
    wire [47:0] _y124;
    wire [47:0] _y125;
    wire [47:0] _y126;
    wire [47:0] _y127;
    GND _gnd (
        .G(gnd)
    );
    VCC _vcc (
        .P(vcc)
    );
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y0 (
        .A({gnd, gnd, gnd, gnd, b0_3[7], b0_3[6], b0_3[5], b0_3[4], b0_3[3], b0_3[2], b0_3[1], b0_3[0], gnd, gnd, gnd, gnd, b0_2[7], b0_2[6], b0_2[5], b0_2[4], b0_2[3], b0_2[2], b0_2[1], b0_2[0], gnd, gnd, gnd, gnd, b0_1[7], b0_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b0_1[5], b0_1[4], b0_1[3], b0_1[2], b0_1[1], b0_1[0], gnd, gnd, gnd, gnd, b0_0[7], b0_0[6], b0_0[5], b0_0[4], b0_0[3], b0_0[2], b0_0[1], b0_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a0_3[7], a0_3[6], a0_3[5], a0_3[4], a0_3[3], a0_3[2], a0_3[1], a0_3[0], gnd, gnd, gnd, gnd, a0_2[7], a0_2[6], a0_2[5], a0_2[4], a0_2[3], a0_2[2], a0_2[1], a0_2[0], gnd, gnd, gnd, gnd, a0_1[7], a0_1[6], a0_1[5], a0_1[4], a0_1[3], a0_1[2], a0_1[1], a0_1[0], gnd, gnd, gnd, gnd, a0_0[7], a0_0[6], a0_0[5], a0_0[4], a0_0[3], a0_0[2], a0_0[1], a0_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y0),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y0_0 = _y0[7:0];
    assign y0_1 = _y0[19:12];
    assign y0_2 = _y0[31:24];
    assign y0_3 = _y0[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y1 (
        .A({gnd, gnd, gnd, gnd, b1_3[7], b1_3[6], b1_3[5], b1_3[4], b1_3[3], b1_3[2], b1_3[1], b1_3[0], gnd, gnd, gnd, gnd, b1_2[7], b1_2[6], b1_2[5], b1_2[4], b1_2[3], b1_2[2], b1_2[1], b1_2[0], gnd, gnd, gnd, gnd, b1_1[7], b1_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b1_1[5], b1_1[4], b1_1[3], b1_1[2], b1_1[1], b1_1[0], gnd, gnd, gnd, gnd, b1_0[7], b1_0[6], b1_0[5], b1_0[4], b1_0[3], b1_0[2], b1_0[1], b1_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a1_3[7], a1_3[6], a1_3[5], a1_3[4], a1_3[3], a1_3[2], a1_3[1], a1_3[0], gnd, gnd, gnd, gnd, a1_2[7], a1_2[6], a1_2[5], a1_2[4], a1_2[3], a1_2[2], a1_2[1], a1_2[0], gnd, gnd, gnd, gnd, a1_1[7], a1_1[6], a1_1[5], a1_1[4], a1_1[3], a1_1[2], a1_1[1], a1_1[0], gnd, gnd, gnd, gnd, a1_0[7], a1_0[6], a1_0[5], a1_0[4], a1_0[3], a1_0[2], a1_0[1], a1_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y1),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y1_0 = _y1[7:0];
    assign y1_1 = _y1[19:12];
    assign y1_2 = _y1[31:24];
    assign y1_3 = _y1[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y2 (
        .A({gnd, gnd, gnd, gnd, b2_3[7], b2_3[6], b2_3[5], b2_3[4], b2_3[3], b2_3[2], b2_3[1], b2_3[0], gnd, gnd, gnd, gnd, b2_2[7], b2_2[6], b2_2[5], b2_2[4], b2_2[3], b2_2[2], b2_2[1], b2_2[0], gnd, gnd, gnd, gnd, b2_1[7], b2_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b2_1[5], b2_1[4], b2_1[3], b2_1[2], b2_1[1], b2_1[0], gnd, gnd, gnd, gnd, b2_0[7], b2_0[6], b2_0[5], b2_0[4], b2_0[3], b2_0[2], b2_0[1], b2_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a2_3[7], a2_3[6], a2_3[5], a2_3[4], a2_3[3], a2_3[2], a2_3[1], a2_3[0], gnd, gnd, gnd, gnd, a2_2[7], a2_2[6], a2_2[5], a2_2[4], a2_2[3], a2_2[2], a2_2[1], a2_2[0], gnd, gnd, gnd, gnd, a2_1[7], a2_1[6], a2_1[5], a2_1[4], a2_1[3], a2_1[2], a2_1[1], a2_1[0], gnd, gnd, gnd, gnd, a2_0[7], a2_0[6], a2_0[5], a2_0[4], a2_0[3], a2_0[2], a2_0[1], a2_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y2),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y2_0 = _y2[7:0];
    assign y2_1 = _y2[19:12];
    assign y2_2 = _y2[31:24];
    assign y2_3 = _y2[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y3 (
        .A({gnd, gnd, gnd, gnd, b3_3[7], b3_3[6], b3_3[5], b3_3[4], b3_3[3], b3_3[2], b3_3[1], b3_3[0], gnd, gnd, gnd, gnd, b3_2[7], b3_2[6], b3_2[5], b3_2[4], b3_2[3], b3_2[2], b3_2[1], b3_2[0], gnd, gnd, gnd, gnd, b3_1[7], b3_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b3_1[5], b3_1[4], b3_1[3], b3_1[2], b3_1[1], b3_1[0], gnd, gnd, gnd, gnd, b3_0[7], b3_0[6], b3_0[5], b3_0[4], b3_0[3], b3_0[2], b3_0[1], b3_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a3_3[7], a3_3[6], a3_3[5], a3_3[4], a3_3[3], a3_3[2], a3_3[1], a3_3[0], gnd, gnd, gnd, gnd, a3_2[7], a3_2[6], a3_2[5], a3_2[4], a3_2[3], a3_2[2], a3_2[1], a3_2[0], gnd, gnd, gnd, gnd, a3_1[7], a3_1[6], a3_1[5], a3_1[4], a3_1[3], a3_1[2], a3_1[1], a3_1[0], gnd, gnd, gnd, gnd, a3_0[7], a3_0[6], a3_0[5], a3_0[4], a3_0[3], a3_0[2], a3_0[1], a3_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y3),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y3_0 = _y3[7:0];
    assign y3_1 = _y3[19:12];
    assign y3_2 = _y3[31:24];
    assign y3_3 = _y3[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y4 (
        .A({gnd, gnd, gnd, gnd, b4_3[7], b4_3[6], b4_3[5], b4_3[4], b4_3[3], b4_3[2], b4_3[1], b4_3[0], gnd, gnd, gnd, gnd, b4_2[7], b4_2[6], b4_2[5], b4_2[4], b4_2[3], b4_2[2], b4_2[1], b4_2[0], gnd, gnd, gnd, gnd, b4_1[7], b4_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b4_1[5], b4_1[4], b4_1[3], b4_1[2], b4_1[1], b4_1[0], gnd, gnd, gnd, gnd, b4_0[7], b4_0[6], b4_0[5], b4_0[4], b4_0[3], b4_0[2], b4_0[1], b4_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a4_3[7], a4_3[6], a4_3[5], a4_3[4], a4_3[3], a4_3[2], a4_3[1], a4_3[0], gnd, gnd, gnd, gnd, a4_2[7], a4_2[6], a4_2[5], a4_2[4], a4_2[3], a4_2[2], a4_2[1], a4_2[0], gnd, gnd, gnd, gnd, a4_1[7], a4_1[6], a4_1[5], a4_1[4], a4_1[3], a4_1[2], a4_1[1], a4_1[0], gnd, gnd, gnd, gnd, a4_0[7], a4_0[6], a4_0[5], a4_0[4], a4_0[3], a4_0[2], a4_0[1], a4_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y4),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y4_0 = _y4[7:0];
    assign y4_1 = _y4[19:12];
    assign y4_2 = _y4[31:24];
    assign y4_3 = _y4[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y5 (
        .A({gnd, gnd, gnd, gnd, b5_3[7], b5_3[6], b5_3[5], b5_3[4], b5_3[3], b5_3[2], b5_3[1], b5_3[0], gnd, gnd, gnd, gnd, b5_2[7], b5_2[6], b5_2[5], b5_2[4], b5_2[3], b5_2[2], b5_2[1], b5_2[0], gnd, gnd, gnd, gnd, b5_1[7], b5_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b5_1[5], b5_1[4], b5_1[3], b5_1[2], b5_1[1], b5_1[0], gnd, gnd, gnd, gnd, b5_0[7], b5_0[6], b5_0[5], b5_0[4], b5_0[3], b5_0[2], b5_0[1], b5_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a5_3[7], a5_3[6], a5_3[5], a5_3[4], a5_3[3], a5_3[2], a5_3[1], a5_3[0], gnd, gnd, gnd, gnd, a5_2[7], a5_2[6], a5_2[5], a5_2[4], a5_2[3], a5_2[2], a5_2[1], a5_2[0], gnd, gnd, gnd, gnd, a5_1[7], a5_1[6], a5_1[5], a5_1[4], a5_1[3], a5_1[2], a5_1[1], a5_1[0], gnd, gnd, gnd, gnd, a5_0[7], a5_0[6], a5_0[5], a5_0[4], a5_0[3], a5_0[2], a5_0[1], a5_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y5),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y5_0 = _y5[7:0];
    assign y5_1 = _y5[19:12];
    assign y5_2 = _y5[31:24];
    assign y5_3 = _y5[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y6 (
        .A({gnd, gnd, gnd, gnd, b6_3[7], b6_3[6], b6_3[5], b6_3[4], b6_3[3], b6_3[2], b6_3[1], b6_3[0], gnd, gnd, gnd, gnd, b6_2[7], b6_2[6], b6_2[5], b6_2[4], b6_2[3], b6_2[2], b6_2[1], b6_2[0], gnd, gnd, gnd, gnd, b6_1[7], b6_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b6_1[5], b6_1[4], b6_1[3], b6_1[2], b6_1[1], b6_1[0], gnd, gnd, gnd, gnd, b6_0[7], b6_0[6], b6_0[5], b6_0[4], b6_0[3], b6_0[2], b6_0[1], b6_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a6_3[7], a6_3[6], a6_3[5], a6_3[4], a6_3[3], a6_3[2], a6_3[1], a6_3[0], gnd, gnd, gnd, gnd, a6_2[7], a6_2[6], a6_2[5], a6_2[4], a6_2[3], a6_2[2], a6_2[1], a6_2[0], gnd, gnd, gnd, gnd, a6_1[7], a6_1[6], a6_1[5], a6_1[4], a6_1[3], a6_1[2], a6_1[1], a6_1[0], gnd, gnd, gnd, gnd, a6_0[7], a6_0[6], a6_0[5], a6_0[4], a6_0[3], a6_0[2], a6_0[1], a6_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y6),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y6_0 = _y6[7:0];
    assign y6_1 = _y6[19:12];
    assign y6_2 = _y6[31:24];
    assign y6_3 = _y6[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y7 (
        .A({gnd, gnd, gnd, gnd, b7_3[7], b7_3[6], b7_3[5], b7_3[4], b7_3[3], b7_3[2], b7_3[1], b7_3[0], gnd, gnd, gnd, gnd, b7_2[7], b7_2[6], b7_2[5], b7_2[4], b7_2[3], b7_2[2], b7_2[1], b7_2[0], gnd, gnd, gnd, gnd, b7_1[7], b7_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b7_1[5], b7_1[4], b7_1[3], b7_1[2], b7_1[1], b7_1[0], gnd, gnd, gnd, gnd, b7_0[7], b7_0[6], b7_0[5], b7_0[4], b7_0[3], b7_0[2], b7_0[1], b7_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a7_3[7], a7_3[6], a7_3[5], a7_3[4], a7_3[3], a7_3[2], a7_3[1], a7_3[0], gnd, gnd, gnd, gnd, a7_2[7], a7_2[6], a7_2[5], a7_2[4], a7_2[3], a7_2[2], a7_2[1], a7_2[0], gnd, gnd, gnd, gnd, a7_1[7], a7_1[6], a7_1[5], a7_1[4], a7_1[3], a7_1[2], a7_1[1], a7_1[0], gnd, gnd, gnd, gnd, a7_0[7], a7_0[6], a7_0[5], a7_0[4], a7_0[3], a7_0[2], a7_0[1], a7_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y7),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y7_0 = _y7[7:0];
    assign y7_1 = _y7[19:12];
    assign y7_2 = _y7[31:24];
    assign y7_3 = _y7[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y8 (
        .A({gnd, gnd, gnd, gnd, b8_3[7], b8_3[6], b8_3[5], b8_3[4], b8_3[3], b8_3[2], b8_3[1], b8_3[0], gnd, gnd, gnd, gnd, b8_2[7], b8_2[6], b8_2[5], b8_2[4], b8_2[3], b8_2[2], b8_2[1], b8_2[0], gnd, gnd, gnd, gnd, b8_1[7], b8_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b8_1[5], b8_1[4], b8_1[3], b8_1[2], b8_1[1], b8_1[0], gnd, gnd, gnd, gnd, b8_0[7], b8_0[6], b8_0[5], b8_0[4], b8_0[3], b8_0[2], b8_0[1], b8_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a8_3[7], a8_3[6], a8_3[5], a8_3[4], a8_3[3], a8_3[2], a8_3[1], a8_3[0], gnd, gnd, gnd, gnd, a8_2[7], a8_2[6], a8_2[5], a8_2[4], a8_2[3], a8_2[2], a8_2[1], a8_2[0], gnd, gnd, gnd, gnd, a8_1[7], a8_1[6], a8_1[5], a8_1[4], a8_1[3], a8_1[2], a8_1[1], a8_1[0], gnd, gnd, gnd, gnd, a8_0[7], a8_0[6], a8_0[5], a8_0[4], a8_0[3], a8_0[2], a8_0[1], a8_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y8),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y8_0 = _y8[7:0];
    assign y8_1 = _y8[19:12];
    assign y8_2 = _y8[31:24];
    assign y8_3 = _y8[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y9 (
        .A({gnd, gnd, gnd, gnd, b9_3[7], b9_3[6], b9_3[5], b9_3[4], b9_3[3], b9_3[2], b9_3[1], b9_3[0], gnd, gnd, gnd, gnd, b9_2[7], b9_2[6], b9_2[5], b9_2[4], b9_2[3], b9_2[2], b9_2[1], b9_2[0], gnd, gnd, gnd, gnd, b9_1[7], b9_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b9_1[5], b9_1[4], b9_1[3], b9_1[2], b9_1[1], b9_1[0], gnd, gnd, gnd, gnd, b9_0[7], b9_0[6], b9_0[5], b9_0[4], b9_0[3], b9_0[2], b9_0[1], b9_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a9_3[7], a9_3[6], a9_3[5], a9_3[4], a9_3[3], a9_3[2], a9_3[1], a9_3[0], gnd, gnd, gnd, gnd, a9_2[7], a9_2[6], a9_2[5], a9_2[4], a9_2[3], a9_2[2], a9_2[1], a9_2[0], gnd, gnd, gnd, gnd, a9_1[7], a9_1[6], a9_1[5], a9_1[4], a9_1[3], a9_1[2], a9_1[1], a9_1[0], gnd, gnd, gnd, gnd, a9_0[7], a9_0[6], a9_0[5], a9_0[4], a9_0[3], a9_0[2], a9_0[1], a9_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y9),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y9_0 = _y9[7:0];
    assign y9_1 = _y9[19:12];
    assign y9_2 = _y9[31:24];
    assign y9_3 = _y9[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y10 (
        .A({gnd, gnd, gnd, gnd, b10_3[7], b10_3[6], b10_3[5], b10_3[4], b10_3[3], b10_3[2], b10_3[1], b10_3[0], gnd, gnd, gnd, gnd, b10_2[7], b10_2[6], b10_2[5], b10_2[4], b10_2[3], b10_2[2], b10_2[1], b10_2[0], gnd, gnd, gnd, gnd, b10_1[7], b10_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b10_1[5], b10_1[4], b10_1[3], b10_1[2], b10_1[1], b10_1[0], gnd, gnd, gnd, gnd, b10_0[7], b10_0[6], b10_0[5], b10_0[4], b10_0[3], b10_0[2], b10_0[1], b10_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a10_3[7], a10_3[6], a10_3[5], a10_3[4], a10_3[3], a10_3[2], a10_3[1], a10_3[0], gnd, gnd, gnd, gnd, a10_2[7], a10_2[6], a10_2[5], a10_2[4], a10_2[3], a10_2[2], a10_2[1], a10_2[0], gnd, gnd, gnd, gnd, a10_1[7], a10_1[6], a10_1[5], a10_1[4], a10_1[3], a10_1[2], a10_1[1], a10_1[0], gnd, gnd, gnd, gnd, a10_0[7], a10_0[6], a10_0[5], a10_0[4], a10_0[3], a10_0[2], a10_0[1], a10_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y10),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y10_0 = _y10[7:0];
    assign y10_1 = _y10[19:12];
    assign y10_2 = _y10[31:24];
    assign y10_3 = _y10[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y11 (
        .A({gnd, gnd, gnd, gnd, b11_3[7], b11_3[6], b11_3[5], b11_3[4], b11_3[3], b11_3[2], b11_3[1], b11_3[0], gnd, gnd, gnd, gnd, b11_2[7], b11_2[6], b11_2[5], b11_2[4], b11_2[3], b11_2[2], b11_2[1], b11_2[0], gnd, gnd, gnd, gnd, b11_1[7], b11_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b11_1[5], b11_1[4], b11_1[3], b11_1[2], b11_1[1], b11_1[0], gnd, gnd, gnd, gnd, b11_0[7], b11_0[6], b11_0[5], b11_0[4], b11_0[3], b11_0[2], b11_0[1], b11_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a11_3[7], a11_3[6], a11_3[5], a11_3[4], a11_3[3], a11_3[2], a11_3[1], a11_3[0], gnd, gnd, gnd, gnd, a11_2[7], a11_2[6], a11_2[5], a11_2[4], a11_2[3], a11_2[2], a11_2[1], a11_2[0], gnd, gnd, gnd, gnd, a11_1[7], a11_1[6], a11_1[5], a11_1[4], a11_1[3], a11_1[2], a11_1[1], a11_1[0], gnd, gnd, gnd, gnd, a11_0[7], a11_0[6], a11_0[5], a11_0[4], a11_0[3], a11_0[2], a11_0[1], a11_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y11),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y11_0 = _y11[7:0];
    assign y11_1 = _y11[19:12];
    assign y11_2 = _y11[31:24];
    assign y11_3 = _y11[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y12 (
        .A({gnd, gnd, gnd, gnd, b12_3[7], b12_3[6], b12_3[5], b12_3[4], b12_3[3], b12_3[2], b12_3[1], b12_3[0], gnd, gnd, gnd, gnd, b12_2[7], b12_2[6], b12_2[5], b12_2[4], b12_2[3], b12_2[2], b12_2[1], b12_2[0], gnd, gnd, gnd, gnd, b12_1[7], b12_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b12_1[5], b12_1[4], b12_1[3], b12_1[2], b12_1[1], b12_1[0], gnd, gnd, gnd, gnd, b12_0[7], b12_0[6], b12_0[5], b12_0[4], b12_0[3], b12_0[2], b12_0[1], b12_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a12_3[7], a12_3[6], a12_3[5], a12_3[4], a12_3[3], a12_3[2], a12_3[1], a12_3[0], gnd, gnd, gnd, gnd, a12_2[7], a12_2[6], a12_2[5], a12_2[4], a12_2[3], a12_2[2], a12_2[1], a12_2[0], gnd, gnd, gnd, gnd, a12_1[7], a12_1[6], a12_1[5], a12_1[4], a12_1[3], a12_1[2], a12_1[1], a12_1[0], gnd, gnd, gnd, gnd, a12_0[7], a12_0[6], a12_0[5], a12_0[4], a12_0[3], a12_0[2], a12_0[1], a12_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y12),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y12_0 = _y12[7:0];
    assign y12_1 = _y12[19:12];
    assign y12_2 = _y12[31:24];
    assign y12_3 = _y12[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y13 (
        .A({gnd, gnd, gnd, gnd, b13_3[7], b13_3[6], b13_3[5], b13_3[4], b13_3[3], b13_3[2], b13_3[1], b13_3[0], gnd, gnd, gnd, gnd, b13_2[7], b13_2[6], b13_2[5], b13_2[4], b13_2[3], b13_2[2], b13_2[1], b13_2[0], gnd, gnd, gnd, gnd, b13_1[7], b13_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b13_1[5], b13_1[4], b13_1[3], b13_1[2], b13_1[1], b13_1[0], gnd, gnd, gnd, gnd, b13_0[7], b13_0[6], b13_0[5], b13_0[4], b13_0[3], b13_0[2], b13_0[1], b13_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a13_3[7], a13_3[6], a13_3[5], a13_3[4], a13_3[3], a13_3[2], a13_3[1], a13_3[0], gnd, gnd, gnd, gnd, a13_2[7], a13_2[6], a13_2[5], a13_2[4], a13_2[3], a13_2[2], a13_2[1], a13_2[0], gnd, gnd, gnd, gnd, a13_1[7], a13_1[6], a13_1[5], a13_1[4], a13_1[3], a13_1[2], a13_1[1], a13_1[0], gnd, gnd, gnd, gnd, a13_0[7], a13_0[6], a13_0[5], a13_0[4], a13_0[3], a13_0[2], a13_0[1], a13_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y13),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y13_0 = _y13[7:0];
    assign y13_1 = _y13[19:12];
    assign y13_2 = _y13[31:24];
    assign y13_3 = _y13[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y14 (
        .A({gnd, gnd, gnd, gnd, b14_3[7], b14_3[6], b14_3[5], b14_3[4], b14_3[3], b14_3[2], b14_3[1], b14_3[0], gnd, gnd, gnd, gnd, b14_2[7], b14_2[6], b14_2[5], b14_2[4], b14_2[3], b14_2[2], b14_2[1], b14_2[0], gnd, gnd, gnd, gnd, b14_1[7], b14_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b14_1[5], b14_1[4], b14_1[3], b14_1[2], b14_1[1], b14_1[0], gnd, gnd, gnd, gnd, b14_0[7], b14_0[6], b14_0[5], b14_0[4], b14_0[3], b14_0[2], b14_0[1], b14_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a14_3[7], a14_3[6], a14_3[5], a14_3[4], a14_3[3], a14_3[2], a14_3[1], a14_3[0], gnd, gnd, gnd, gnd, a14_2[7], a14_2[6], a14_2[5], a14_2[4], a14_2[3], a14_2[2], a14_2[1], a14_2[0], gnd, gnd, gnd, gnd, a14_1[7], a14_1[6], a14_1[5], a14_1[4], a14_1[3], a14_1[2], a14_1[1], a14_1[0], gnd, gnd, gnd, gnd, a14_0[7], a14_0[6], a14_0[5], a14_0[4], a14_0[3], a14_0[2], a14_0[1], a14_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y14),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y14_0 = _y14[7:0];
    assign y14_1 = _y14[19:12];
    assign y14_2 = _y14[31:24];
    assign y14_3 = _y14[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y15 (
        .A({gnd, gnd, gnd, gnd, b15_3[7], b15_3[6], b15_3[5], b15_3[4], b15_3[3], b15_3[2], b15_3[1], b15_3[0], gnd, gnd, gnd, gnd, b15_2[7], b15_2[6], b15_2[5], b15_2[4], b15_2[3], b15_2[2], b15_2[1], b15_2[0], gnd, gnd, gnd, gnd, b15_1[7], b15_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b15_1[5], b15_1[4], b15_1[3], b15_1[2], b15_1[1], b15_1[0], gnd, gnd, gnd, gnd, b15_0[7], b15_0[6], b15_0[5], b15_0[4], b15_0[3], b15_0[2], b15_0[1], b15_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a15_3[7], a15_3[6], a15_3[5], a15_3[4], a15_3[3], a15_3[2], a15_3[1], a15_3[0], gnd, gnd, gnd, gnd, a15_2[7], a15_2[6], a15_2[5], a15_2[4], a15_2[3], a15_2[2], a15_2[1], a15_2[0], gnd, gnd, gnd, gnd, a15_1[7], a15_1[6], a15_1[5], a15_1[4], a15_1[3], a15_1[2], a15_1[1], a15_1[0], gnd, gnd, gnd, gnd, a15_0[7], a15_0[6], a15_0[5], a15_0[4], a15_0[3], a15_0[2], a15_0[1], a15_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y15),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y15_0 = _y15[7:0];
    assign y15_1 = _y15[19:12];
    assign y15_2 = _y15[31:24];
    assign y15_3 = _y15[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y16 (
        .A({gnd, gnd, gnd, gnd, b16_3[7], b16_3[6], b16_3[5], b16_3[4], b16_3[3], b16_3[2], b16_3[1], b16_3[0], gnd, gnd, gnd, gnd, b16_2[7], b16_2[6], b16_2[5], b16_2[4], b16_2[3], b16_2[2], b16_2[1], b16_2[0], gnd, gnd, gnd, gnd, b16_1[7], b16_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b16_1[5], b16_1[4], b16_1[3], b16_1[2], b16_1[1], b16_1[0], gnd, gnd, gnd, gnd, b16_0[7], b16_0[6], b16_0[5], b16_0[4], b16_0[3], b16_0[2], b16_0[1], b16_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a16_3[7], a16_3[6], a16_3[5], a16_3[4], a16_3[3], a16_3[2], a16_3[1], a16_3[0], gnd, gnd, gnd, gnd, a16_2[7], a16_2[6], a16_2[5], a16_2[4], a16_2[3], a16_2[2], a16_2[1], a16_2[0], gnd, gnd, gnd, gnd, a16_1[7], a16_1[6], a16_1[5], a16_1[4], a16_1[3], a16_1[2], a16_1[1], a16_1[0], gnd, gnd, gnd, gnd, a16_0[7], a16_0[6], a16_0[5], a16_0[4], a16_0[3], a16_0[2], a16_0[1], a16_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y16),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y16_0 = _y16[7:0];
    assign y16_1 = _y16[19:12];
    assign y16_2 = _y16[31:24];
    assign y16_3 = _y16[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y17 (
        .A({gnd, gnd, gnd, gnd, b17_3[7], b17_3[6], b17_3[5], b17_3[4], b17_3[3], b17_3[2], b17_3[1], b17_3[0], gnd, gnd, gnd, gnd, b17_2[7], b17_2[6], b17_2[5], b17_2[4], b17_2[3], b17_2[2], b17_2[1], b17_2[0], gnd, gnd, gnd, gnd, b17_1[7], b17_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b17_1[5], b17_1[4], b17_1[3], b17_1[2], b17_1[1], b17_1[0], gnd, gnd, gnd, gnd, b17_0[7], b17_0[6], b17_0[5], b17_0[4], b17_0[3], b17_0[2], b17_0[1], b17_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a17_3[7], a17_3[6], a17_3[5], a17_3[4], a17_3[3], a17_3[2], a17_3[1], a17_3[0], gnd, gnd, gnd, gnd, a17_2[7], a17_2[6], a17_2[5], a17_2[4], a17_2[3], a17_2[2], a17_2[1], a17_2[0], gnd, gnd, gnd, gnd, a17_1[7], a17_1[6], a17_1[5], a17_1[4], a17_1[3], a17_1[2], a17_1[1], a17_1[0], gnd, gnd, gnd, gnd, a17_0[7], a17_0[6], a17_0[5], a17_0[4], a17_0[3], a17_0[2], a17_0[1], a17_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y17),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y17_0 = _y17[7:0];
    assign y17_1 = _y17[19:12];
    assign y17_2 = _y17[31:24];
    assign y17_3 = _y17[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y18 (
        .A({gnd, gnd, gnd, gnd, b18_3[7], b18_3[6], b18_3[5], b18_3[4], b18_3[3], b18_3[2], b18_3[1], b18_3[0], gnd, gnd, gnd, gnd, b18_2[7], b18_2[6], b18_2[5], b18_2[4], b18_2[3], b18_2[2], b18_2[1], b18_2[0], gnd, gnd, gnd, gnd, b18_1[7], b18_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b18_1[5], b18_1[4], b18_1[3], b18_1[2], b18_1[1], b18_1[0], gnd, gnd, gnd, gnd, b18_0[7], b18_0[6], b18_0[5], b18_0[4], b18_0[3], b18_0[2], b18_0[1], b18_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a18_3[7], a18_3[6], a18_3[5], a18_3[4], a18_3[3], a18_3[2], a18_3[1], a18_3[0], gnd, gnd, gnd, gnd, a18_2[7], a18_2[6], a18_2[5], a18_2[4], a18_2[3], a18_2[2], a18_2[1], a18_2[0], gnd, gnd, gnd, gnd, a18_1[7], a18_1[6], a18_1[5], a18_1[4], a18_1[3], a18_1[2], a18_1[1], a18_1[0], gnd, gnd, gnd, gnd, a18_0[7], a18_0[6], a18_0[5], a18_0[4], a18_0[3], a18_0[2], a18_0[1], a18_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y18),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y18_0 = _y18[7:0];
    assign y18_1 = _y18[19:12];
    assign y18_2 = _y18[31:24];
    assign y18_3 = _y18[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y19 (
        .A({gnd, gnd, gnd, gnd, b19_3[7], b19_3[6], b19_3[5], b19_3[4], b19_3[3], b19_3[2], b19_3[1], b19_3[0], gnd, gnd, gnd, gnd, b19_2[7], b19_2[6], b19_2[5], b19_2[4], b19_2[3], b19_2[2], b19_2[1], b19_2[0], gnd, gnd, gnd, gnd, b19_1[7], b19_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b19_1[5], b19_1[4], b19_1[3], b19_1[2], b19_1[1], b19_1[0], gnd, gnd, gnd, gnd, b19_0[7], b19_0[6], b19_0[5], b19_0[4], b19_0[3], b19_0[2], b19_0[1], b19_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a19_3[7], a19_3[6], a19_3[5], a19_3[4], a19_3[3], a19_3[2], a19_3[1], a19_3[0], gnd, gnd, gnd, gnd, a19_2[7], a19_2[6], a19_2[5], a19_2[4], a19_2[3], a19_2[2], a19_2[1], a19_2[0], gnd, gnd, gnd, gnd, a19_1[7], a19_1[6], a19_1[5], a19_1[4], a19_1[3], a19_1[2], a19_1[1], a19_1[0], gnd, gnd, gnd, gnd, a19_0[7], a19_0[6], a19_0[5], a19_0[4], a19_0[3], a19_0[2], a19_0[1], a19_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y19),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y19_0 = _y19[7:0];
    assign y19_1 = _y19[19:12];
    assign y19_2 = _y19[31:24];
    assign y19_3 = _y19[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y20 (
        .A({gnd, gnd, gnd, gnd, b20_3[7], b20_3[6], b20_3[5], b20_3[4], b20_3[3], b20_3[2], b20_3[1], b20_3[0], gnd, gnd, gnd, gnd, b20_2[7], b20_2[6], b20_2[5], b20_2[4], b20_2[3], b20_2[2], b20_2[1], b20_2[0], gnd, gnd, gnd, gnd, b20_1[7], b20_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b20_1[5], b20_1[4], b20_1[3], b20_1[2], b20_1[1], b20_1[0], gnd, gnd, gnd, gnd, b20_0[7], b20_0[6], b20_0[5], b20_0[4], b20_0[3], b20_0[2], b20_0[1], b20_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a20_3[7], a20_3[6], a20_3[5], a20_3[4], a20_3[3], a20_3[2], a20_3[1], a20_3[0], gnd, gnd, gnd, gnd, a20_2[7], a20_2[6], a20_2[5], a20_2[4], a20_2[3], a20_2[2], a20_2[1], a20_2[0], gnd, gnd, gnd, gnd, a20_1[7], a20_1[6], a20_1[5], a20_1[4], a20_1[3], a20_1[2], a20_1[1], a20_1[0], gnd, gnd, gnd, gnd, a20_0[7], a20_0[6], a20_0[5], a20_0[4], a20_0[3], a20_0[2], a20_0[1], a20_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y20),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y20_0 = _y20[7:0];
    assign y20_1 = _y20[19:12];
    assign y20_2 = _y20[31:24];
    assign y20_3 = _y20[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y21 (
        .A({gnd, gnd, gnd, gnd, b21_3[7], b21_3[6], b21_3[5], b21_3[4], b21_3[3], b21_3[2], b21_3[1], b21_3[0], gnd, gnd, gnd, gnd, b21_2[7], b21_2[6], b21_2[5], b21_2[4], b21_2[3], b21_2[2], b21_2[1], b21_2[0], gnd, gnd, gnd, gnd, b21_1[7], b21_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b21_1[5], b21_1[4], b21_1[3], b21_1[2], b21_1[1], b21_1[0], gnd, gnd, gnd, gnd, b21_0[7], b21_0[6], b21_0[5], b21_0[4], b21_0[3], b21_0[2], b21_0[1], b21_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a21_3[7], a21_3[6], a21_3[5], a21_3[4], a21_3[3], a21_3[2], a21_3[1], a21_3[0], gnd, gnd, gnd, gnd, a21_2[7], a21_2[6], a21_2[5], a21_2[4], a21_2[3], a21_2[2], a21_2[1], a21_2[0], gnd, gnd, gnd, gnd, a21_1[7], a21_1[6], a21_1[5], a21_1[4], a21_1[3], a21_1[2], a21_1[1], a21_1[0], gnd, gnd, gnd, gnd, a21_0[7], a21_0[6], a21_0[5], a21_0[4], a21_0[3], a21_0[2], a21_0[1], a21_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y21),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y21_0 = _y21[7:0];
    assign y21_1 = _y21[19:12];
    assign y21_2 = _y21[31:24];
    assign y21_3 = _y21[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y22 (
        .A({gnd, gnd, gnd, gnd, b22_3[7], b22_3[6], b22_3[5], b22_3[4], b22_3[3], b22_3[2], b22_3[1], b22_3[0], gnd, gnd, gnd, gnd, b22_2[7], b22_2[6], b22_2[5], b22_2[4], b22_2[3], b22_2[2], b22_2[1], b22_2[0], gnd, gnd, gnd, gnd, b22_1[7], b22_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b22_1[5], b22_1[4], b22_1[3], b22_1[2], b22_1[1], b22_1[0], gnd, gnd, gnd, gnd, b22_0[7], b22_0[6], b22_0[5], b22_0[4], b22_0[3], b22_0[2], b22_0[1], b22_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a22_3[7], a22_3[6], a22_3[5], a22_3[4], a22_3[3], a22_3[2], a22_3[1], a22_3[0], gnd, gnd, gnd, gnd, a22_2[7], a22_2[6], a22_2[5], a22_2[4], a22_2[3], a22_2[2], a22_2[1], a22_2[0], gnd, gnd, gnd, gnd, a22_1[7], a22_1[6], a22_1[5], a22_1[4], a22_1[3], a22_1[2], a22_1[1], a22_1[0], gnd, gnd, gnd, gnd, a22_0[7], a22_0[6], a22_0[5], a22_0[4], a22_0[3], a22_0[2], a22_0[1], a22_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y22),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y22_0 = _y22[7:0];
    assign y22_1 = _y22[19:12];
    assign y22_2 = _y22[31:24];
    assign y22_3 = _y22[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y23 (
        .A({gnd, gnd, gnd, gnd, b23_3[7], b23_3[6], b23_3[5], b23_3[4], b23_3[3], b23_3[2], b23_3[1], b23_3[0], gnd, gnd, gnd, gnd, b23_2[7], b23_2[6], b23_2[5], b23_2[4], b23_2[3], b23_2[2], b23_2[1], b23_2[0], gnd, gnd, gnd, gnd, b23_1[7], b23_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b23_1[5], b23_1[4], b23_1[3], b23_1[2], b23_1[1], b23_1[0], gnd, gnd, gnd, gnd, b23_0[7], b23_0[6], b23_0[5], b23_0[4], b23_0[3], b23_0[2], b23_0[1], b23_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a23_3[7], a23_3[6], a23_3[5], a23_3[4], a23_3[3], a23_3[2], a23_3[1], a23_3[0], gnd, gnd, gnd, gnd, a23_2[7], a23_2[6], a23_2[5], a23_2[4], a23_2[3], a23_2[2], a23_2[1], a23_2[0], gnd, gnd, gnd, gnd, a23_1[7], a23_1[6], a23_1[5], a23_1[4], a23_1[3], a23_1[2], a23_1[1], a23_1[0], gnd, gnd, gnd, gnd, a23_0[7], a23_0[6], a23_0[5], a23_0[4], a23_0[3], a23_0[2], a23_0[1], a23_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y23),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y23_0 = _y23[7:0];
    assign y23_1 = _y23[19:12];
    assign y23_2 = _y23[31:24];
    assign y23_3 = _y23[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y24 (
        .A({gnd, gnd, gnd, gnd, b24_3[7], b24_3[6], b24_3[5], b24_3[4], b24_3[3], b24_3[2], b24_3[1], b24_3[0], gnd, gnd, gnd, gnd, b24_2[7], b24_2[6], b24_2[5], b24_2[4], b24_2[3], b24_2[2], b24_2[1], b24_2[0], gnd, gnd, gnd, gnd, b24_1[7], b24_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b24_1[5], b24_1[4], b24_1[3], b24_1[2], b24_1[1], b24_1[0], gnd, gnd, gnd, gnd, b24_0[7], b24_0[6], b24_0[5], b24_0[4], b24_0[3], b24_0[2], b24_0[1], b24_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a24_3[7], a24_3[6], a24_3[5], a24_3[4], a24_3[3], a24_3[2], a24_3[1], a24_3[0], gnd, gnd, gnd, gnd, a24_2[7], a24_2[6], a24_2[5], a24_2[4], a24_2[3], a24_2[2], a24_2[1], a24_2[0], gnd, gnd, gnd, gnd, a24_1[7], a24_1[6], a24_1[5], a24_1[4], a24_1[3], a24_1[2], a24_1[1], a24_1[0], gnd, gnd, gnd, gnd, a24_0[7], a24_0[6], a24_0[5], a24_0[4], a24_0[3], a24_0[2], a24_0[1], a24_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y24),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y24_0 = _y24[7:0];
    assign y24_1 = _y24[19:12];
    assign y24_2 = _y24[31:24];
    assign y24_3 = _y24[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y25 (
        .A({gnd, gnd, gnd, gnd, b25_3[7], b25_3[6], b25_3[5], b25_3[4], b25_3[3], b25_3[2], b25_3[1], b25_3[0], gnd, gnd, gnd, gnd, b25_2[7], b25_2[6], b25_2[5], b25_2[4], b25_2[3], b25_2[2], b25_2[1], b25_2[0], gnd, gnd, gnd, gnd, b25_1[7], b25_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b25_1[5], b25_1[4], b25_1[3], b25_1[2], b25_1[1], b25_1[0], gnd, gnd, gnd, gnd, b25_0[7], b25_0[6], b25_0[5], b25_0[4], b25_0[3], b25_0[2], b25_0[1], b25_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a25_3[7], a25_3[6], a25_3[5], a25_3[4], a25_3[3], a25_3[2], a25_3[1], a25_3[0], gnd, gnd, gnd, gnd, a25_2[7], a25_2[6], a25_2[5], a25_2[4], a25_2[3], a25_2[2], a25_2[1], a25_2[0], gnd, gnd, gnd, gnd, a25_1[7], a25_1[6], a25_1[5], a25_1[4], a25_1[3], a25_1[2], a25_1[1], a25_1[0], gnd, gnd, gnd, gnd, a25_0[7], a25_0[6], a25_0[5], a25_0[4], a25_0[3], a25_0[2], a25_0[1], a25_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y25),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y25_0 = _y25[7:0];
    assign y25_1 = _y25[19:12];
    assign y25_2 = _y25[31:24];
    assign y25_3 = _y25[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y26 (
        .A({gnd, gnd, gnd, gnd, b26_3[7], b26_3[6], b26_3[5], b26_3[4], b26_3[3], b26_3[2], b26_3[1], b26_3[0], gnd, gnd, gnd, gnd, b26_2[7], b26_2[6], b26_2[5], b26_2[4], b26_2[3], b26_2[2], b26_2[1], b26_2[0], gnd, gnd, gnd, gnd, b26_1[7], b26_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b26_1[5], b26_1[4], b26_1[3], b26_1[2], b26_1[1], b26_1[0], gnd, gnd, gnd, gnd, b26_0[7], b26_0[6], b26_0[5], b26_0[4], b26_0[3], b26_0[2], b26_0[1], b26_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a26_3[7], a26_3[6], a26_3[5], a26_3[4], a26_3[3], a26_3[2], a26_3[1], a26_3[0], gnd, gnd, gnd, gnd, a26_2[7], a26_2[6], a26_2[5], a26_2[4], a26_2[3], a26_2[2], a26_2[1], a26_2[0], gnd, gnd, gnd, gnd, a26_1[7], a26_1[6], a26_1[5], a26_1[4], a26_1[3], a26_1[2], a26_1[1], a26_1[0], gnd, gnd, gnd, gnd, a26_0[7], a26_0[6], a26_0[5], a26_0[4], a26_0[3], a26_0[2], a26_0[1], a26_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y26),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y26_0 = _y26[7:0];
    assign y26_1 = _y26[19:12];
    assign y26_2 = _y26[31:24];
    assign y26_3 = _y26[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y27 (
        .A({gnd, gnd, gnd, gnd, b27_3[7], b27_3[6], b27_3[5], b27_3[4], b27_3[3], b27_3[2], b27_3[1], b27_3[0], gnd, gnd, gnd, gnd, b27_2[7], b27_2[6], b27_2[5], b27_2[4], b27_2[3], b27_2[2], b27_2[1], b27_2[0], gnd, gnd, gnd, gnd, b27_1[7], b27_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b27_1[5], b27_1[4], b27_1[3], b27_1[2], b27_1[1], b27_1[0], gnd, gnd, gnd, gnd, b27_0[7], b27_0[6], b27_0[5], b27_0[4], b27_0[3], b27_0[2], b27_0[1], b27_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a27_3[7], a27_3[6], a27_3[5], a27_3[4], a27_3[3], a27_3[2], a27_3[1], a27_3[0], gnd, gnd, gnd, gnd, a27_2[7], a27_2[6], a27_2[5], a27_2[4], a27_2[3], a27_2[2], a27_2[1], a27_2[0], gnd, gnd, gnd, gnd, a27_1[7], a27_1[6], a27_1[5], a27_1[4], a27_1[3], a27_1[2], a27_1[1], a27_1[0], gnd, gnd, gnd, gnd, a27_0[7], a27_0[6], a27_0[5], a27_0[4], a27_0[3], a27_0[2], a27_0[1], a27_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y27),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y27_0 = _y27[7:0];
    assign y27_1 = _y27[19:12];
    assign y27_2 = _y27[31:24];
    assign y27_3 = _y27[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y28 (
        .A({gnd, gnd, gnd, gnd, b28_3[7], b28_3[6], b28_3[5], b28_3[4], b28_3[3], b28_3[2], b28_3[1], b28_3[0], gnd, gnd, gnd, gnd, b28_2[7], b28_2[6], b28_2[5], b28_2[4], b28_2[3], b28_2[2], b28_2[1], b28_2[0], gnd, gnd, gnd, gnd, b28_1[7], b28_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b28_1[5], b28_1[4], b28_1[3], b28_1[2], b28_1[1], b28_1[0], gnd, gnd, gnd, gnd, b28_0[7], b28_0[6], b28_0[5], b28_0[4], b28_0[3], b28_0[2], b28_0[1], b28_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a28_3[7], a28_3[6], a28_3[5], a28_3[4], a28_3[3], a28_3[2], a28_3[1], a28_3[0], gnd, gnd, gnd, gnd, a28_2[7], a28_2[6], a28_2[5], a28_2[4], a28_2[3], a28_2[2], a28_2[1], a28_2[0], gnd, gnd, gnd, gnd, a28_1[7], a28_1[6], a28_1[5], a28_1[4], a28_1[3], a28_1[2], a28_1[1], a28_1[0], gnd, gnd, gnd, gnd, a28_0[7], a28_0[6], a28_0[5], a28_0[4], a28_0[3], a28_0[2], a28_0[1], a28_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y28),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y28_0 = _y28[7:0];
    assign y28_1 = _y28[19:12];
    assign y28_2 = _y28[31:24];
    assign y28_3 = _y28[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y29 (
        .A({gnd, gnd, gnd, gnd, b29_3[7], b29_3[6], b29_3[5], b29_3[4], b29_3[3], b29_3[2], b29_3[1], b29_3[0], gnd, gnd, gnd, gnd, b29_2[7], b29_2[6], b29_2[5], b29_2[4], b29_2[3], b29_2[2], b29_2[1], b29_2[0], gnd, gnd, gnd, gnd, b29_1[7], b29_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b29_1[5], b29_1[4], b29_1[3], b29_1[2], b29_1[1], b29_1[0], gnd, gnd, gnd, gnd, b29_0[7], b29_0[6], b29_0[5], b29_0[4], b29_0[3], b29_0[2], b29_0[1], b29_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a29_3[7], a29_3[6], a29_3[5], a29_3[4], a29_3[3], a29_3[2], a29_3[1], a29_3[0], gnd, gnd, gnd, gnd, a29_2[7], a29_2[6], a29_2[5], a29_2[4], a29_2[3], a29_2[2], a29_2[1], a29_2[0], gnd, gnd, gnd, gnd, a29_1[7], a29_1[6], a29_1[5], a29_1[4], a29_1[3], a29_1[2], a29_1[1], a29_1[0], gnd, gnd, gnd, gnd, a29_0[7], a29_0[6], a29_0[5], a29_0[4], a29_0[3], a29_0[2], a29_0[1], a29_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y29),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y29_0 = _y29[7:0];
    assign y29_1 = _y29[19:12];
    assign y29_2 = _y29[31:24];
    assign y29_3 = _y29[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y30 (
        .A({gnd, gnd, gnd, gnd, b30_3[7], b30_3[6], b30_3[5], b30_3[4], b30_3[3], b30_3[2], b30_3[1], b30_3[0], gnd, gnd, gnd, gnd, b30_2[7], b30_2[6], b30_2[5], b30_2[4], b30_2[3], b30_2[2], b30_2[1], b30_2[0], gnd, gnd, gnd, gnd, b30_1[7], b30_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b30_1[5], b30_1[4], b30_1[3], b30_1[2], b30_1[1], b30_1[0], gnd, gnd, gnd, gnd, b30_0[7], b30_0[6], b30_0[5], b30_0[4], b30_0[3], b30_0[2], b30_0[1], b30_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a30_3[7], a30_3[6], a30_3[5], a30_3[4], a30_3[3], a30_3[2], a30_3[1], a30_3[0], gnd, gnd, gnd, gnd, a30_2[7], a30_2[6], a30_2[5], a30_2[4], a30_2[3], a30_2[2], a30_2[1], a30_2[0], gnd, gnd, gnd, gnd, a30_1[7], a30_1[6], a30_1[5], a30_1[4], a30_1[3], a30_1[2], a30_1[1], a30_1[0], gnd, gnd, gnd, gnd, a30_0[7], a30_0[6], a30_0[5], a30_0[4], a30_0[3], a30_0[2], a30_0[1], a30_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y30),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y30_0 = _y30[7:0];
    assign y30_1 = _y30[19:12];
    assign y30_2 = _y30[31:24];
    assign y30_3 = _y30[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y31 (
        .A({gnd, gnd, gnd, gnd, b31_3[7], b31_3[6], b31_3[5], b31_3[4], b31_3[3], b31_3[2], b31_3[1], b31_3[0], gnd, gnd, gnd, gnd, b31_2[7], b31_2[6], b31_2[5], b31_2[4], b31_2[3], b31_2[2], b31_2[1], b31_2[0], gnd, gnd, gnd, gnd, b31_1[7], b31_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b31_1[5], b31_1[4], b31_1[3], b31_1[2], b31_1[1], b31_1[0], gnd, gnd, gnd, gnd, b31_0[7], b31_0[6], b31_0[5], b31_0[4], b31_0[3], b31_0[2], b31_0[1], b31_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a31_3[7], a31_3[6], a31_3[5], a31_3[4], a31_3[3], a31_3[2], a31_3[1], a31_3[0], gnd, gnd, gnd, gnd, a31_2[7], a31_2[6], a31_2[5], a31_2[4], a31_2[3], a31_2[2], a31_2[1], a31_2[0], gnd, gnd, gnd, gnd, a31_1[7], a31_1[6], a31_1[5], a31_1[4], a31_1[3], a31_1[2], a31_1[1], a31_1[0], gnd, gnd, gnd, gnd, a31_0[7], a31_0[6], a31_0[5], a31_0[4], a31_0[3], a31_0[2], a31_0[1], a31_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y31),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y31_0 = _y31[7:0];
    assign y31_1 = _y31[19:12];
    assign y31_2 = _y31[31:24];
    assign y31_3 = _y31[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y32 (
        .A({gnd, gnd, gnd, gnd, b32_3[7], b32_3[6], b32_3[5], b32_3[4], b32_3[3], b32_3[2], b32_3[1], b32_3[0], gnd, gnd, gnd, gnd, b32_2[7], b32_2[6], b32_2[5], b32_2[4], b32_2[3], b32_2[2], b32_2[1], b32_2[0], gnd, gnd, gnd, gnd, b32_1[7], b32_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b32_1[5], b32_1[4], b32_1[3], b32_1[2], b32_1[1], b32_1[0], gnd, gnd, gnd, gnd, b32_0[7], b32_0[6], b32_0[5], b32_0[4], b32_0[3], b32_0[2], b32_0[1], b32_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a32_3[7], a32_3[6], a32_3[5], a32_3[4], a32_3[3], a32_3[2], a32_3[1], a32_3[0], gnd, gnd, gnd, gnd, a32_2[7], a32_2[6], a32_2[5], a32_2[4], a32_2[3], a32_2[2], a32_2[1], a32_2[0], gnd, gnd, gnd, gnd, a32_1[7], a32_1[6], a32_1[5], a32_1[4], a32_1[3], a32_1[2], a32_1[1], a32_1[0], gnd, gnd, gnd, gnd, a32_0[7], a32_0[6], a32_0[5], a32_0[4], a32_0[3], a32_0[2], a32_0[1], a32_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y32),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y32_0 = _y32[7:0];
    assign y32_1 = _y32[19:12];
    assign y32_2 = _y32[31:24];
    assign y32_3 = _y32[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y33 (
        .A({gnd, gnd, gnd, gnd, b33_3[7], b33_3[6], b33_3[5], b33_3[4], b33_3[3], b33_3[2], b33_3[1], b33_3[0], gnd, gnd, gnd, gnd, b33_2[7], b33_2[6], b33_2[5], b33_2[4], b33_2[3], b33_2[2], b33_2[1], b33_2[0], gnd, gnd, gnd, gnd, b33_1[7], b33_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b33_1[5], b33_1[4], b33_1[3], b33_1[2], b33_1[1], b33_1[0], gnd, gnd, gnd, gnd, b33_0[7], b33_0[6], b33_0[5], b33_0[4], b33_0[3], b33_0[2], b33_0[1], b33_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a33_3[7], a33_3[6], a33_3[5], a33_3[4], a33_3[3], a33_3[2], a33_3[1], a33_3[0], gnd, gnd, gnd, gnd, a33_2[7], a33_2[6], a33_2[5], a33_2[4], a33_2[3], a33_2[2], a33_2[1], a33_2[0], gnd, gnd, gnd, gnd, a33_1[7], a33_1[6], a33_1[5], a33_1[4], a33_1[3], a33_1[2], a33_1[1], a33_1[0], gnd, gnd, gnd, gnd, a33_0[7], a33_0[6], a33_0[5], a33_0[4], a33_0[3], a33_0[2], a33_0[1], a33_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y33),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y33_0 = _y33[7:0];
    assign y33_1 = _y33[19:12];
    assign y33_2 = _y33[31:24];
    assign y33_3 = _y33[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y34 (
        .A({gnd, gnd, gnd, gnd, b34_3[7], b34_3[6], b34_3[5], b34_3[4], b34_3[3], b34_3[2], b34_3[1], b34_3[0], gnd, gnd, gnd, gnd, b34_2[7], b34_2[6], b34_2[5], b34_2[4], b34_2[3], b34_2[2], b34_2[1], b34_2[0], gnd, gnd, gnd, gnd, b34_1[7], b34_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b34_1[5], b34_1[4], b34_1[3], b34_1[2], b34_1[1], b34_1[0], gnd, gnd, gnd, gnd, b34_0[7], b34_0[6], b34_0[5], b34_0[4], b34_0[3], b34_0[2], b34_0[1], b34_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a34_3[7], a34_3[6], a34_3[5], a34_3[4], a34_3[3], a34_3[2], a34_3[1], a34_3[0], gnd, gnd, gnd, gnd, a34_2[7], a34_2[6], a34_2[5], a34_2[4], a34_2[3], a34_2[2], a34_2[1], a34_2[0], gnd, gnd, gnd, gnd, a34_1[7], a34_1[6], a34_1[5], a34_1[4], a34_1[3], a34_1[2], a34_1[1], a34_1[0], gnd, gnd, gnd, gnd, a34_0[7], a34_0[6], a34_0[5], a34_0[4], a34_0[3], a34_0[2], a34_0[1], a34_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y34),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y34_0 = _y34[7:0];
    assign y34_1 = _y34[19:12];
    assign y34_2 = _y34[31:24];
    assign y34_3 = _y34[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y35 (
        .A({gnd, gnd, gnd, gnd, b35_3[7], b35_3[6], b35_3[5], b35_3[4], b35_3[3], b35_3[2], b35_3[1], b35_3[0], gnd, gnd, gnd, gnd, b35_2[7], b35_2[6], b35_2[5], b35_2[4], b35_2[3], b35_2[2], b35_2[1], b35_2[0], gnd, gnd, gnd, gnd, b35_1[7], b35_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b35_1[5], b35_1[4], b35_1[3], b35_1[2], b35_1[1], b35_1[0], gnd, gnd, gnd, gnd, b35_0[7], b35_0[6], b35_0[5], b35_0[4], b35_0[3], b35_0[2], b35_0[1], b35_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a35_3[7], a35_3[6], a35_3[5], a35_3[4], a35_3[3], a35_3[2], a35_3[1], a35_3[0], gnd, gnd, gnd, gnd, a35_2[7], a35_2[6], a35_2[5], a35_2[4], a35_2[3], a35_2[2], a35_2[1], a35_2[0], gnd, gnd, gnd, gnd, a35_1[7], a35_1[6], a35_1[5], a35_1[4], a35_1[3], a35_1[2], a35_1[1], a35_1[0], gnd, gnd, gnd, gnd, a35_0[7], a35_0[6], a35_0[5], a35_0[4], a35_0[3], a35_0[2], a35_0[1], a35_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y35),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y35_0 = _y35[7:0];
    assign y35_1 = _y35[19:12];
    assign y35_2 = _y35[31:24];
    assign y35_3 = _y35[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y36 (
        .A({gnd, gnd, gnd, gnd, b36_3[7], b36_3[6], b36_3[5], b36_3[4], b36_3[3], b36_3[2], b36_3[1], b36_3[0], gnd, gnd, gnd, gnd, b36_2[7], b36_2[6], b36_2[5], b36_2[4], b36_2[3], b36_2[2], b36_2[1], b36_2[0], gnd, gnd, gnd, gnd, b36_1[7], b36_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b36_1[5], b36_1[4], b36_1[3], b36_1[2], b36_1[1], b36_1[0], gnd, gnd, gnd, gnd, b36_0[7], b36_0[6], b36_0[5], b36_0[4], b36_0[3], b36_0[2], b36_0[1], b36_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a36_3[7], a36_3[6], a36_3[5], a36_3[4], a36_3[3], a36_3[2], a36_3[1], a36_3[0], gnd, gnd, gnd, gnd, a36_2[7], a36_2[6], a36_2[5], a36_2[4], a36_2[3], a36_2[2], a36_2[1], a36_2[0], gnd, gnd, gnd, gnd, a36_1[7], a36_1[6], a36_1[5], a36_1[4], a36_1[3], a36_1[2], a36_1[1], a36_1[0], gnd, gnd, gnd, gnd, a36_0[7], a36_0[6], a36_0[5], a36_0[4], a36_0[3], a36_0[2], a36_0[1], a36_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y36),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y36_0 = _y36[7:0];
    assign y36_1 = _y36[19:12];
    assign y36_2 = _y36[31:24];
    assign y36_3 = _y36[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y37 (
        .A({gnd, gnd, gnd, gnd, b37_3[7], b37_3[6], b37_3[5], b37_3[4], b37_3[3], b37_3[2], b37_3[1], b37_3[0], gnd, gnd, gnd, gnd, b37_2[7], b37_2[6], b37_2[5], b37_2[4], b37_2[3], b37_2[2], b37_2[1], b37_2[0], gnd, gnd, gnd, gnd, b37_1[7], b37_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b37_1[5], b37_1[4], b37_1[3], b37_1[2], b37_1[1], b37_1[0], gnd, gnd, gnd, gnd, b37_0[7], b37_0[6], b37_0[5], b37_0[4], b37_0[3], b37_0[2], b37_0[1], b37_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a37_3[7], a37_3[6], a37_3[5], a37_3[4], a37_3[3], a37_3[2], a37_3[1], a37_3[0], gnd, gnd, gnd, gnd, a37_2[7], a37_2[6], a37_2[5], a37_2[4], a37_2[3], a37_2[2], a37_2[1], a37_2[0], gnd, gnd, gnd, gnd, a37_1[7], a37_1[6], a37_1[5], a37_1[4], a37_1[3], a37_1[2], a37_1[1], a37_1[0], gnd, gnd, gnd, gnd, a37_0[7], a37_0[6], a37_0[5], a37_0[4], a37_0[3], a37_0[2], a37_0[1], a37_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y37),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y37_0 = _y37[7:0];
    assign y37_1 = _y37[19:12];
    assign y37_2 = _y37[31:24];
    assign y37_3 = _y37[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y38 (
        .A({gnd, gnd, gnd, gnd, b38_3[7], b38_3[6], b38_3[5], b38_3[4], b38_3[3], b38_3[2], b38_3[1], b38_3[0], gnd, gnd, gnd, gnd, b38_2[7], b38_2[6], b38_2[5], b38_2[4], b38_2[3], b38_2[2], b38_2[1], b38_2[0], gnd, gnd, gnd, gnd, b38_1[7], b38_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b38_1[5], b38_1[4], b38_1[3], b38_1[2], b38_1[1], b38_1[0], gnd, gnd, gnd, gnd, b38_0[7], b38_0[6], b38_0[5], b38_0[4], b38_0[3], b38_0[2], b38_0[1], b38_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a38_3[7], a38_3[6], a38_3[5], a38_3[4], a38_3[3], a38_3[2], a38_3[1], a38_3[0], gnd, gnd, gnd, gnd, a38_2[7], a38_2[6], a38_2[5], a38_2[4], a38_2[3], a38_2[2], a38_2[1], a38_2[0], gnd, gnd, gnd, gnd, a38_1[7], a38_1[6], a38_1[5], a38_1[4], a38_1[3], a38_1[2], a38_1[1], a38_1[0], gnd, gnd, gnd, gnd, a38_0[7], a38_0[6], a38_0[5], a38_0[4], a38_0[3], a38_0[2], a38_0[1], a38_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y38),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y38_0 = _y38[7:0];
    assign y38_1 = _y38[19:12];
    assign y38_2 = _y38[31:24];
    assign y38_3 = _y38[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y39 (
        .A({gnd, gnd, gnd, gnd, b39_3[7], b39_3[6], b39_3[5], b39_3[4], b39_3[3], b39_3[2], b39_3[1], b39_3[0], gnd, gnd, gnd, gnd, b39_2[7], b39_2[6], b39_2[5], b39_2[4], b39_2[3], b39_2[2], b39_2[1], b39_2[0], gnd, gnd, gnd, gnd, b39_1[7], b39_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b39_1[5], b39_1[4], b39_1[3], b39_1[2], b39_1[1], b39_1[0], gnd, gnd, gnd, gnd, b39_0[7], b39_0[6], b39_0[5], b39_0[4], b39_0[3], b39_0[2], b39_0[1], b39_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a39_3[7], a39_3[6], a39_3[5], a39_3[4], a39_3[3], a39_3[2], a39_3[1], a39_3[0], gnd, gnd, gnd, gnd, a39_2[7], a39_2[6], a39_2[5], a39_2[4], a39_2[3], a39_2[2], a39_2[1], a39_2[0], gnd, gnd, gnd, gnd, a39_1[7], a39_1[6], a39_1[5], a39_1[4], a39_1[3], a39_1[2], a39_1[1], a39_1[0], gnd, gnd, gnd, gnd, a39_0[7], a39_0[6], a39_0[5], a39_0[4], a39_0[3], a39_0[2], a39_0[1], a39_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y39),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y39_0 = _y39[7:0];
    assign y39_1 = _y39[19:12];
    assign y39_2 = _y39[31:24];
    assign y39_3 = _y39[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y40 (
        .A({gnd, gnd, gnd, gnd, b40_3[7], b40_3[6], b40_3[5], b40_3[4], b40_3[3], b40_3[2], b40_3[1], b40_3[0], gnd, gnd, gnd, gnd, b40_2[7], b40_2[6], b40_2[5], b40_2[4], b40_2[3], b40_2[2], b40_2[1], b40_2[0], gnd, gnd, gnd, gnd, b40_1[7], b40_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b40_1[5], b40_1[4], b40_1[3], b40_1[2], b40_1[1], b40_1[0], gnd, gnd, gnd, gnd, b40_0[7], b40_0[6], b40_0[5], b40_0[4], b40_0[3], b40_0[2], b40_0[1], b40_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a40_3[7], a40_3[6], a40_3[5], a40_3[4], a40_3[3], a40_3[2], a40_3[1], a40_3[0], gnd, gnd, gnd, gnd, a40_2[7], a40_2[6], a40_2[5], a40_2[4], a40_2[3], a40_2[2], a40_2[1], a40_2[0], gnd, gnd, gnd, gnd, a40_1[7], a40_1[6], a40_1[5], a40_1[4], a40_1[3], a40_1[2], a40_1[1], a40_1[0], gnd, gnd, gnd, gnd, a40_0[7], a40_0[6], a40_0[5], a40_0[4], a40_0[3], a40_0[2], a40_0[1], a40_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y40),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y40_0 = _y40[7:0];
    assign y40_1 = _y40[19:12];
    assign y40_2 = _y40[31:24];
    assign y40_3 = _y40[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y41 (
        .A({gnd, gnd, gnd, gnd, b41_3[7], b41_3[6], b41_3[5], b41_3[4], b41_3[3], b41_3[2], b41_3[1], b41_3[0], gnd, gnd, gnd, gnd, b41_2[7], b41_2[6], b41_2[5], b41_2[4], b41_2[3], b41_2[2], b41_2[1], b41_2[0], gnd, gnd, gnd, gnd, b41_1[7], b41_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b41_1[5], b41_1[4], b41_1[3], b41_1[2], b41_1[1], b41_1[0], gnd, gnd, gnd, gnd, b41_0[7], b41_0[6], b41_0[5], b41_0[4], b41_0[3], b41_0[2], b41_0[1], b41_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a41_3[7], a41_3[6], a41_3[5], a41_3[4], a41_3[3], a41_3[2], a41_3[1], a41_3[0], gnd, gnd, gnd, gnd, a41_2[7], a41_2[6], a41_2[5], a41_2[4], a41_2[3], a41_2[2], a41_2[1], a41_2[0], gnd, gnd, gnd, gnd, a41_1[7], a41_1[6], a41_1[5], a41_1[4], a41_1[3], a41_1[2], a41_1[1], a41_1[0], gnd, gnd, gnd, gnd, a41_0[7], a41_0[6], a41_0[5], a41_0[4], a41_0[3], a41_0[2], a41_0[1], a41_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y41),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y41_0 = _y41[7:0];
    assign y41_1 = _y41[19:12];
    assign y41_2 = _y41[31:24];
    assign y41_3 = _y41[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y42 (
        .A({gnd, gnd, gnd, gnd, b42_3[7], b42_3[6], b42_3[5], b42_3[4], b42_3[3], b42_3[2], b42_3[1], b42_3[0], gnd, gnd, gnd, gnd, b42_2[7], b42_2[6], b42_2[5], b42_2[4], b42_2[3], b42_2[2], b42_2[1], b42_2[0], gnd, gnd, gnd, gnd, b42_1[7], b42_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b42_1[5], b42_1[4], b42_1[3], b42_1[2], b42_1[1], b42_1[0], gnd, gnd, gnd, gnd, b42_0[7], b42_0[6], b42_0[5], b42_0[4], b42_0[3], b42_0[2], b42_0[1], b42_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a42_3[7], a42_3[6], a42_3[5], a42_3[4], a42_3[3], a42_3[2], a42_3[1], a42_3[0], gnd, gnd, gnd, gnd, a42_2[7], a42_2[6], a42_2[5], a42_2[4], a42_2[3], a42_2[2], a42_2[1], a42_2[0], gnd, gnd, gnd, gnd, a42_1[7], a42_1[6], a42_1[5], a42_1[4], a42_1[3], a42_1[2], a42_1[1], a42_1[0], gnd, gnd, gnd, gnd, a42_0[7], a42_0[6], a42_0[5], a42_0[4], a42_0[3], a42_0[2], a42_0[1], a42_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y42),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y42_0 = _y42[7:0];
    assign y42_1 = _y42[19:12];
    assign y42_2 = _y42[31:24];
    assign y42_3 = _y42[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y43 (
        .A({gnd, gnd, gnd, gnd, b43_3[7], b43_3[6], b43_3[5], b43_3[4], b43_3[3], b43_3[2], b43_3[1], b43_3[0], gnd, gnd, gnd, gnd, b43_2[7], b43_2[6], b43_2[5], b43_2[4], b43_2[3], b43_2[2], b43_2[1], b43_2[0], gnd, gnd, gnd, gnd, b43_1[7], b43_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b43_1[5], b43_1[4], b43_1[3], b43_1[2], b43_1[1], b43_1[0], gnd, gnd, gnd, gnd, b43_0[7], b43_0[6], b43_0[5], b43_0[4], b43_0[3], b43_0[2], b43_0[1], b43_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a43_3[7], a43_3[6], a43_3[5], a43_3[4], a43_3[3], a43_3[2], a43_3[1], a43_3[0], gnd, gnd, gnd, gnd, a43_2[7], a43_2[6], a43_2[5], a43_2[4], a43_2[3], a43_2[2], a43_2[1], a43_2[0], gnd, gnd, gnd, gnd, a43_1[7], a43_1[6], a43_1[5], a43_1[4], a43_1[3], a43_1[2], a43_1[1], a43_1[0], gnd, gnd, gnd, gnd, a43_0[7], a43_0[6], a43_0[5], a43_0[4], a43_0[3], a43_0[2], a43_0[1], a43_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y43),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y43_0 = _y43[7:0];
    assign y43_1 = _y43[19:12];
    assign y43_2 = _y43[31:24];
    assign y43_3 = _y43[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y44 (
        .A({gnd, gnd, gnd, gnd, b44_3[7], b44_3[6], b44_3[5], b44_3[4], b44_3[3], b44_3[2], b44_3[1], b44_3[0], gnd, gnd, gnd, gnd, b44_2[7], b44_2[6], b44_2[5], b44_2[4], b44_2[3], b44_2[2], b44_2[1], b44_2[0], gnd, gnd, gnd, gnd, b44_1[7], b44_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b44_1[5], b44_1[4], b44_1[3], b44_1[2], b44_1[1], b44_1[0], gnd, gnd, gnd, gnd, b44_0[7], b44_0[6], b44_0[5], b44_0[4], b44_0[3], b44_0[2], b44_0[1], b44_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a44_3[7], a44_3[6], a44_3[5], a44_3[4], a44_3[3], a44_3[2], a44_3[1], a44_3[0], gnd, gnd, gnd, gnd, a44_2[7], a44_2[6], a44_2[5], a44_2[4], a44_2[3], a44_2[2], a44_2[1], a44_2[0], gnd, gnd, gnd, gnd, a44_1[7], a44_1[6], a44_1[5], a44_1[4], a44_1[3], a44_1[2], a44_1[1], a44_1[0], gnd, gnd, gnd, gnd, a44_0[7], a44_0[6], a44_0[5], a44_0[4], a44_0[3], a44_0[2], a44_0[1], a44_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y44),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y44_0 = _y44[7:0];
    assign y44_1 = _y44[19:12];
    assign y44_2 = _y44[31:24];
    assign y44_3 = _y44[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y45 (
        .A({gnd, gnd, gnd, gnd, b45_3[7], b45_3[6], b45_3[5], b45_3[4], b45_3[3], b45_3[2], b45_3[1], b45_3[0], gnd, gnd, gnd, gnd, b45_2[7], b45_2[6], b45_2[5], b45_2[4], b45_2[3], b45_2[2], b45_2[1], b45_2[0], gnd, gnd, gnd, gnd, b45_1[7], b45_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b45_1[5], b45_1[4], b45_1[3], b45_1[2], b45_1[1], b45_1[0], gnd, gnd, gnd, gnd, b45_0[7], b45_0[6], b45_0[5], b45_0[4], b45_0[3], b45_0[2], b45_0[1], b45_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a45_3[7], a45_3[6], a45_3[5], a45_3[4], a45_3[3], a45_3[2], a45_3[1], a45_3[0], gnd, gnd, gnd, gnd, a45_2[7], a45_2[6], a45_2[5], a45_2[4], a45_2[3], a45_2[2], a45_2[1], a45_2[0], gnd, gnd, gnd, gnd, a45_1[7], a45_1[6], a45_1[5], a45_1[4], a45_1[3], a45_1[2], a45_1[1], a45_1[0], gnd, gnd, gnd, gnd, a45_0[7], a45_0[6], a45_0[5], a45_0[4], a45_0[3], a45_0[2], a45_0[1], a45_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y45),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y45_0 = _y45[7:0];
    assign y45_1 = _y45[19:12];
    assign y45_2 = _y45[31:24];
    assign y45_3 = _y45[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y46 (
        .A({gnd, gnd, gnd, gnd, b46_3[7], b46_3[6], b46_3[5], b46_3[4], b46_3[3], b46_3[2], b46_3[1], b46_3[0], gnd, gnd, gnd, gnd, b46_2[7], b46_2[6], b46_2[5], b46_2[4], b46_2[3], b46_2[2], b46_2[1], b46_2[0], gnd, gnd, gnd, gnd, b46_1[7], b46_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b46_1[5], b46_1[4], b46_1[3], b46_1[2], b46_1[1], b46_1[0], gnd, gnd, gnd, gnd, b46_0[7], b46_0[6], b46_0[5], b46_0[4], b46_0[3], b46_0[2], b46_0[1], b46_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a46_3[7], a46_3[6], a46_3[5], a46_3[4], a46_3[3], a46_3[2], a46_3[1], a46_3[0], gnd, gnd, gnd, gnd, a46_2[7], a46_2[6], a46_2[5], a46_2[4], a46_2[3], a46_2[2], a46_2[1], a46_2[0], gnd, gnd, gnd, gnd, a46_1[7], a46_1[6], a46_1[5], a46_1[4], a46_1[3], a46_1[2], a46_1[1], a46_1[0], gnd, gnd, gnd, gnd, a46_0[7], a46_0[6], a46_0[5], a46_0[4], a46_0[3], a46_0[2], a46_0[1], a46_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y46),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y46_0 = _y46[7:0];
    assign y46_1 = _y46[19:12];
    assign y46_2 = _y46[31:24];
    assign y46_3 = _y46[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y47 (
        .A({gnd, gnd, gnd, gnd, b47_3[7], b47_3[6], b47_3[5], b47_3[4], b47_3[3], b47_3[2], b47_3[1], b47_3[0], gnd, gnd, gnd, gnd, b47_2[7], b47_2[6], b47_2[5], b47_2[4], b47_2[3], b47_2[2], b47_2[1], b47_2[0], gnd, gnd, gnd, gnd, b47_1[7], b47_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b47_1[5], b47_1[4], b47_1[3], b47_1[2], b47_1[1], b47_1[0], gnd, gnd, gnd, gnd, b47_0[7], b47_0[6], b47_0[5], b47_0[4], b47_0[3], b47_0[2], b47_0[1], b47_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a47_3[7], a47_3[6], a47_3[5], a47_3[4], a47_3[3], a47_3[2], a47_3[1], a47_3[0], gnd, gnd, gnd, gnd, a47_2[7], a47_2[6], a47_2[5], a47_2[4], a47_2[3], a47_2[2], a47_2[1], a47_2[0], gnd, gnd, gnd, gnd, a47_1[7], a47_1[6], a47_1[5], a47_1[4], a47_1[3], a47_1[2], a47_1[1], a47_1[0], gnd, gnd, gnd, gnd, a47_0[7], a47_0[6], a47_0[5], a47_0[4], a47_0[3], a47_0[2], a47_0[1], a47_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y47),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y47_0 = _y47[7:0];
    assign y47_1 = _y47[19:12];
    assign y47_2 = _y47[31:24];
    assign y47_3 = _y47[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y48 (
        .A({gnd, gnd, gnd, gnd, b48_3[7], b48_3[6], b48_3[5], b48_3[4], b48_3[3], b48_3[2], b48_3[1], b48_3[0], gnd, gnd, gnd, gnd, b48_2[7], b48_2[6], b48_2[5], b48_2[4], b48_2[3], b48_2[2], b48_2[1], b48_2[0], gnd, gnd, gnd, gnd, b48_1[7], b48_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b48_1[5], b48_1[4], b48_1[3], b48_1[2], b48_1[1], b48_1[0], gnd, gnd, gnd, gnd, b48_0[7], b48_0[6], b48_0[5], b48_0[4], b48_0[3], b48_0[2], b48_0[1], b48_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a48_3[7], a48_3[6], a48_3[5], a48_3[4], a48_3[3], a48_3[2], a48_3[1], a48_3[0], gnd, gnd, gnd, gnd, a48_2[7], a48_2[6], a48_2[5], a48_2[4], a48_2[3], a48_2[2], a48_2[1], a48_2[0], gnd, gnd, gnd, gnd, a48_1[7], a48_1[6], a48_1[5], a48_1[4], a48_1[3], a48_1[2], a48_1[1], a48_1[0], gnd, gnd, gnd, gnd, a48_0[7], a48_0[6], a48_0[5], a48_0[4], a48_0[3], a48_0[2], a48_0[1], a48_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y48),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y48_0 = _y48[7:0];
    assign y48_1 = _y48[19:12];
    assign y48_2 = _y48[31:24];
    assign y48_3 = _y48[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y49 (
        .A({gnd, gnd, gnd, gnd, b49_3[7], b49_3[6], b49_3[5], b49_3[4], b49_3[3], b49_3[2], b49_3[1], b49_3[0], gnd, gnd, gnd, gnd, b49_2[7], b49_2[6], b49_2[5], b49_2[4], b49_2[3], b49_2[2], b49_2[1], b49_2[0], gnd, gnd, gnd, gnd, b49_1[7], b49_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b49_1[5], b49_1[4], b49_1[3], b49_1[2], b49_1[1], b49_1[0], gnd, gnd, gnd, gnd, b49_0[7], b49_0[6], b49_0[5], b49_0[4], b49_0[3], b49_0[2], b49_0[1], b49_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a49_3[7], a49_3[6], a49_3[5], a49_3[4], a49_3[3], a49_3[2], a49_3[1], a49_3[0], gnd, gnd, gnd, gnd, a49_2[7], a49_2[6], a49_2[5], a49_2[4], a49_2[3], a49_2[2], a49_2[1], a49_2[0], gnd, gnd, gnd, gnd, a49_1[7], a49_1[6], a49_1[5], a49_1[4], a49_1[3], a49_1[2], a49_1[1], a49_1[0], gnd, gnd, gnd, gnd, a49_0[7], a49_0[6], a49_0[5], a49_0[4], a49_0[3], a49_0[2], a49_0[1], a49_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y49),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y49_0 = _y49[7:0];
    assign y49_1 = _y49[19:12];
    assign y49_2 = _y49[31:24];
    assign y49_3 = _y49[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y50 (
        .A({gnd, gnd, gnd, gnd, b50_3[7], b50_3[6], b50_3[5], b50_3[4], b50_3[3], b50_3[2], b50_3[1], b50_3[0], gnd, gnd, gnd, gnd, b50_2[7], b50_2[6], b50_2[5], b50_2[4], b50_2[3], b50_2[2], b50_2[1], b50_2[0], gnd, gnd, gnd, gnd, b50_1[7], b50_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b50_1[5], b50_1[4], b50_1[3], b50_1[2], b50_1[1], b50_1[0], gnd, gnd, gnd, gnd, b50_0[7], b50_0[6], b50_0[5], b50_0[4], b50_0[3], b50_0[2], b50_0[1], b50_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a50_3[7], a50_3[6], a50_3[5], a50_3[4], a50_3[3], a50_3[2], a50_3[1], a50_3[0], gnd, gnd, gnd, gnd, a50_2[7], a50_2[6], a50_2[5], a50_2[4], a50_2[3], a50_2[2], a50_2[1], a50_2[0], gnd, gnd, gnd, gnd, a50_1[7], a50_1[6], a50_1[5], a50_1[4], a50_1[3], a50_1[2], a50_1[1], a50_1[0], gnd, gnd, gnd, gnd, a50_0[7], a50_0[6], a50_0[5], a50_0[4], a50_0[3], a50_0[2], a50_0[1], a50_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y50),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y50_0 = _y50[7:0];
    assign y50_1 = _y50[19:12];
    assign y50_2 = _y50[31:24];
    assign y50_3 = _y50[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y51 (
        .A({gnd, gnd, gnd, gnd, b51_3[7], b51_3[6], b51_3[5], b51_3[4], b51_3[3], b51_3[2], b51_3[1], b51_3[0], gnd, gnd, gnd, gnd, b51_2[7], b51_2[6], b51_2[5], b51_2[4], b51_2[3], b51_2[2], b51_2[1], b51_2[0], gnd, gnd, gnd, gnd, b51_1[7], b51_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b51_1[5], b51_1[4], b51_1[3], b51_1[2], b51_1[1], b51_1[0], gnd, gnd, gnd, gnd, b51_0[7], b51_0[6], b51_0[5], b51_0[4], b51_0[3], b51_0[2], b51_0[1], b51_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a51_3[7], a51_3[6], a51_3[5], a51_3[4], a51_3[3], a51_3[2], a51_3[1], a51_3[0], gnd, gnd, gnd, gnd, a51_2[7], a51_2[6], a51_2[5], a51_2[4], a51_2[3], a51_2[2], a51_2[1], a51_2[0], gnd, gnd, gnd, gnd, a51_1[7], a51_1[6], a51_1[5], a51_1[4], a51_1[3], a51_1[2], a51_1[1], a51_1[0], gnd, gnd, gnd, gnd, a51_0[7], a51_0[6], a51_0[5], a51_0[4], a51_0[3], a51_0[2], a51_0[1], a51_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y51),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y51_0 = _y51[7:0];
    assign y51_1 = _y51[19:12];
    assign y51_2 = _y51[31:24];
    assign y51_3 = _y51[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y52 (
        .A({gnd, gnd, gnd, gnd, b52_3[7], b52_3[6], b52_3[5], b52_3[4], b52_3[3], b52_3[2], b52_3[1], b52_3[0], gnd, gnd, gnd, gnd, b52_2[7], b52_2[6], b52_2[5], b52_2[4], b52_2[3], b52_2[2], b52_2[1], b52_2[0], gnd, gnd, gnd, gnd, b52_1[7], b52_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b52_1[5], b52_1[4], b52_1[3], b52_1[2], b52_1[1], b52_1[0], gnd, gnd, gnd, gnd, b52_0[7], b52_0[6], b52_0[5], b52_0[4], b52_0[3], b52_0[2], b52_0[1], b52_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a52_3[7], a52_3[6], a52_3[5], a52_3[4], a52_3[3], a52_3[2], a52_3[1], a52_3[0], gnd, gnd, gnd, gnd, a52_2[7], a52_2[6], a52_2[5], a52_2[4], a52_2[3], a52_2[2], a52_2[1], a52_2[0], gnd, gnd, gnd, gnd, a52_1[7], a52_1[6], a52_1[5], a52_1[4], a52_1[3], a52_1[2], a52_1[1], a52_1[0], gnd, gnd, gnd, gnd, a52_0[7], a52_0[6], a52_0[5], a52_0[4], a52_0[3], a52_0[2], a52_0[1], a52_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y52),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y52_0 = _y52[7:0];
    assign y52_1 = _y52[19:12];
    assign y52_2 = _y52[31:24];
    assign y52_3 = _y52[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y53 (
        .A({gnd, gnd, gnd, gnd, b53_3[7], b53_3[6], b53_3[5], b53_3[4], b53_3[3], b53_3[2], b53_3[1], b53_3[0], gnd, gnd, gnd, gnd, b53_2[7], b53_2[6], b53_2[5], b53_2[4], b53_2[3], b53_2[2], b53_2[1], b53_2[0], gnd, gnd, gnd, gnd, b53_1[7], b53_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b53_1[5], b53_1[4], b53_1[3], b53_1[2], b53_1[1], b53_1[0], gnd, gnd, gnd, gnd, b53_0[7], b53_0[6], b53_0[5], b53_0[4], b53_0[3], b53_0[2], b53_0[1], b53_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a53_3[7], a53_3[6], a53_3[5], a53_3[4], a53_3[3], a53_3[2], a53_3[1], a53_3[0], gnd, gnd, gnd, gnd, a53_2[7], a53_2[6], a53_2[5], a53_2[4], a53_2[3], a53_2[2], a53_2[1], a53_2[0], gnd, gnd, gnd, gnd, a53_1[7], a53_1[6], a53_1[5], a53_1[4], a53_1[3], a53_1[2], a53_1[1], a53_1[0], gnd, gnd, gnd, gnd, a53_0[7], a53_0[6], a53_0[5], a53_0[4], a53_0[3], a53_0[2], a53_0[1], a53_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y53),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y53_0 = _y53[7:0];
    assign y53_1 = _y53[19:12];
    assign y53_2 = _y53[31:24];
    assign y53_3 = _y53[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y54 (
        .A({gnd, gnd, gnd, gnd, b54_3[7], b54_3[6], b54_3[5], b54_3[4], b54_3[3], b54_3[2], b54_3[1], b54_3[0], gnd, gnd, gnd, gnd, b54_2[7], b54_2[6], b54_2[5], b54_2[4], b54_2[3], b54_2[2], b54_2[1], b54_2[0], gnd, gnd, gnd, gnd, b54_1[7], b54_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b54_1[5], b54_1[4], b54_1[3], b54_1[2], b54_1[1], b54_1[0], gnd, gnd, gnd, gnd, b54_0[7], b54_0[6], b54_0[5], b54_0[4], b54_0[3], b54_0[2], b54_0[1], b54_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a54_3[7], a54_3[6], a54_3[5], a54_3[4], a54_3[3], a54_3[2], a54_3[1], a54_3[0], gnd, gnd, gnd, gnd, a54_2[7], a54_2[6], a54_2[5], a54_2[4], a54_2[3], a54_2[2], a54_2[1], a54_2[0], gnd, gnd, gnd, gnd, a54_1[7], a54_1[6], a54_1[5], a54_1[4], a54_1[3], a54_1[2], a54_1[1], a54_1[0], gnd, gnd, gnd, gnd, a54_0[7], a54_0[6], a54_0[5], a54_0[4], a54_0[3], a54_0[2], a54_0[1], a54_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y54),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y54_0 = _y54[7:0];
    assign y54_1 = _y54[19:12];
    assign y54_2 = _y54[31:24];
    assign y54_3 = _y54[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y55 (
        .A({gnd, gnd, gnd, gnd, b55_3[7], b55_3[6], b55_3[5], b55_3[4], b55_3[3], b55_3[2], b55_3[1], b55_3[0], gnd, gnd, gnd, gnd, b55_2[7], b55_2[6], b55_2[5], b55_2[4], b55_2[3], b55_2[2], b55_2[1], b55_2[0], gnd, gnd, gnd, gnd, b55_1[7], b55_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b55_1[5], b55_1[4], b55_1[3], b55_1[2], b55_1[1], b55_1[0], gnd, gnd, gnd, gnd, b55_0[7], b55_0[6], b55_0[5], b55_0[4], b55_0[3], b55_0[2], b55_0[1], b55_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a55_3[7], a55_3[6], a55_3[5], a55_3[4], a55_3[3], a55_3[2], a55_3[1], a55_3[0], gnd, gnd, gnd, gnd, a55_2[7], a55_2[6], a55_2[5], a55_2[4], a55_2[3], a55_2[2], a55_2[1], a55_2[0], gnd, gnd, gnd, gnd, a55_1[7], a55_1[6], a55_1[5], a55_1[4], a55_1[3], a55_1[2], a55_1[1], a55_1[0], gnd, gnd, gnd, gnd, a55_0[7], a55_0[6], a55_0[5], a55_0[4], a55_0[3], a55_0[2], a55_0[1], a55_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y55),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y55_0 = _y55[7:0];
    assign y55_1 = _y55[19:12];
    assign y55_2 = _y55[31:24];
    assign y55_3 = _y55[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y56 (
        .A({gnd, gnd, gnd, gnd, b56_3[7], b56_3[6], b56_3[5], b56_3[4], b56_3[3], b56_3[2], b56_3[1], b56_3[0], gnd, gnd, gnd, gnd, b56_2[7], b56_2[6], b56_2[5], b56_2[4], b56_2[3], b56_2[2], b56_2[1], b56_2[0], gnd, gnd, gnd, gnd, b56_1[7], b56_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b56_1[5], b56_1[4], b56_1[3], b56_1[2], b56_1[1], b56_1[0], gnd, gnd, gnd, gnd, b56_0[7], b56_0[6], b56_0[5], b56_0[4], b56_0[3], b56_0[2], b56_0[1], b56_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a56_3[7], a56_3[6], a56_3[5], a56_3[4], a56_3[3], a56_3[2], a56_3[1], a56_3[0], gnd, gnd, gnd, gnd, a56_2[7], a56_2[6], a56_2[5], a56_2[4], a56_2[3], a56_2[2], a56_2[1], a56_2[0], gnd, gnd, gnd, gnd, a56_1[7], a56_1[6], a56_1[5], a56_1[4], a56_1[3], a56_1[2], a56_1[1], a56_1[0], gnd, gnd, gnd, gnd, a56_0[7], a56_0[6], a56_0[5], a56_0[4], a56_0[3], a56_0[2], a56_0[1], a56_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y56),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y56_0 = _y56[7:0];
    assign y56_1 = _y56[19:12];
    assign y56_2 = _y56[31:24];
    assign y56_3 = _y56[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y57 (
        .A({gnd, gnd, gnd, gnd, b57_3[7], b57_3[6], b57_3[5], b57_3[4], b57_3[3], b57_3[2], b57_3[1], b57_3[0], gnd, gnd, gnd, gnd, b57_2[7], b57_2[6], b57_2[5], b57_2[4], b57_2[3], b57_2[2], b57_2[1], b57_2[0], gnd, gnd, gnd, gnd, b57_1[7], b57_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b57_1[5], b57_1[4], b57_1[3], b57_1[2], b57_1[1], b57_1[0], gnd, gnd, gnd, gnd, b57_0[7], b57_0[6], b57_0[5], b57_0[4], b57_0[3], b57_0[2], b57_0[1], b57_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a57_3[7], a57_3[6], a57_3[5], a57_3[4], a57_3[3], a57_3[2], a57_3[1], a57_3[0], gnd, gnd, gnd, gnd, a57_2[7], a57_2[6], a57_2[5], a57_2[4], a57_2[3], a57_2[2], a57_2[1], a57_2[0], gnd, gnd, gnd, gnd, a57_1[7], a57_1[6], a57_1[5], a57_1[4], a57_1[3], a57_1[2], a57_1[1], a57_1[0], gnd, gnd, gnd, gnd, a57_0[7], a57_0[6], a57_0[5], a57_0[4], a57_0[3], a57_0[2], a57_0[1], a57_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y57),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y57_0 = _y57[7:0];
    assign y57_1 = _y57[19:12];
    assign y57_2 = _y57[31:24];
    assign y57_3 = _y57[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y58 (
        .A({gnd, gnd, gnd, gnd, b58_3[7], b58_3[6], b58_3[5], b58_3[4], b58_3[3], b58_3[2], b58_3[1], b58_3[0], gnd, gnd, gnd, gnd, b58_2[7], b58_2[6], b58_2[5], b58_2[4], b58_2[3], b58_2[2], b58_2[1], b58_2[0], gnd, gnd, gnd, gnd, b58_1[7], b58_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b58_1[5], b58_1[4], b58_1[3], b58_1[2], b58_1[1], b58_1[0], gnd, gnd, gnd, gnd, b58_0[7], b58_0[6], b58_0[5], b58_0[4], b58_0[3], b58_0[2], b58_0[1], b58_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a58_3[7], a58_3[6], a58_3[5], a58_3[4], a58_3[3], a58_3[2], a58_3[1], a58_3[0], gnd, gnd, gnd, gnd, a58_2[7], a58_2[6], a58_2[5], a58_2[4], a58_2[3], a58_2[2], a58_2[1], a58_2[0], gnd, gnd, gnd, gnd, a58_1[7], a58_1[6], a58_1[5], a58_1[4], a58_1[3], a58_1[2], a58_1[1], a58_1[0], gnd, gnd, gnd, gnd, a58_0[7], a58_0[6], a58_0[5], a58_0[4], a58_0[3], a58_0[2], a58_0[1], a58_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y58),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y58_0 = _y58[7:0];
    assign y58_1 = _y58[19:12];
    assign y58_2 = _y58[31:24];
    assign y58_3 = _y58[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y59 (
        .A({gnd, gnd, gnd, gnd, b59_3[7], b59_3[6], b59_3[5], b59_3[4], b59_3[3], b59_3[2], b59_3[1], b59_3[0], gnd, gnd, gnd, gnd, b59_2[7], b59_2[6], b59_2[5], b59_2[4], b59_2[3], b59_2[2], b59_2[1], b59_2[0], gnd, gnd, gnd, gnd, b59_1[7], b59_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b59_1[5], b59_1[4], b59_1[3], b59_1[2], b59_1[1], b59_1[0], gnd, gnd, gnd, gnd, b59_0[7], b59_0[6], b59_0[5], b59_0[4], b59_0[3], b59_0[2], b59_0[1], b59_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a59_3[7], a59_3[6], a59_3[5], a59_3[4], a59_3[3], a59_3[2], a59_3[1], a59_3[0], gnd, gnd, gnd, gnd, a59_2[7], a59_2[6], a59_2[5], a59_2[4], a59_2[3], a59_2[2], a59_2[1], a59_2[0], gnd, gnd, gnd, gnd, a59_1[7], a59_1[6], a59_1[5], a59_1[4], a59_1[3], a59_1[2], a59_1[1], a59_1[0], gnd, gnd, gnd, gnd, a59_0[7], a59_0[6], a59_0[5], a59_0[4], a59_0[3], a59_0[2], a59_0[1], a59_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y59),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y59_0 = _y59[7:0];
    assign y59_1 = _y59[19:12];
    assign y59_2 = _y59[31:24];
    assign y59_3 = _y59[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y60 (
        .A({gnd, gnd, gnd, gnd, b60_3[7], b60_3[6], b60_3[5], b60_3[4], b60_3[3], b60_3[2], b60_3[1], b60_3[0], gnd, gnd, gnd, gnd, b60_2[7], b60_2[6], b60_2[5], b60_2[4], b60_2[3], b60_2[2], b60_2[1], b60_2[0], gnd, gnd, gnd, gnd, b60_1[7], b60_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b60_1[5], b60_1[4], b60_1[3], b60_1[2], b60_1[1], b60_1[0], gnd, gnd, gnd, gnd, b60_0[7], b60_0[6], b60_0[5], b60_0[4], b60_0[3], b60_0[2], b60_0[1], b60_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a60_3[7], a60_3[6], a60_3[5], a60_3[4], a60_3[3], a60_3[2], a60_3[1], a60_3[0], gnd, gnd, gnd, gnd, a60_2[7], a60_2[6], a60_2[5], a60_2[4], a60_2[3], a60_2[2], a60_2[1], a60_2[0], gnd, gnd, gnd, gnd, a60_1[7], a60_1[6], a60_1[5], a60_1[4], a60_1[3], a60_1[2], a60_1[1], a60_1[0], gnd, gnd, gnd, gnd, a60_0[7], a60_0[6], a60_0[5], a60_0[4], a60_0[3], a60_0[2], a60_0[1], a60_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y60),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y60_0 = _y60[7:0];
    assign y60_1 = _y60[19:12];
    assign y60_2 = _y60[31:24];
    assign y60_3 = _y60[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y61 (
        .A({gnd, gnd, gnd, gnd, b61_3[7], b61_3[6], b61_3[5], b61_3[4], b61_3[3], b61_3[2], b61_3[1], b61_3[0], gnd, gnd, gnd, gnd, b61_2[7], b61_2[6], b61_2[5], b61_2[4], b61_2[3], b61_2[2], b61_2[1], b61_2[0], gnd, gnd, gnd, gnd, b61_1[7], b61_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b61_1[5], b61_1[4], b61_1[3], b61_1[2], b61_1[1], b61_1[0], gnd, gnd, gnd, gnd, b61_0[7], b61_0[6], b61_0[5], b61_0[4], b61_0[3], b61_0[2], b61_0[1], b61_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a61_3[7], a61_3[6], a61_3[5], a61_3[4], a61_3[3], a61_3[2], a61_3[1], a61_3[0], gnd, gnd, gnd, gnd, a61_2[7], a61_2[6], a61_2[5], a61_2[4], a61_2[3], a61_2[2], a61_2[1], a61_2[0], gnd, gnd, gnd, gnd, a61_1[7], a61_1[6], a61_1[5], a61_1[4], a61_1[3], a61_1[2], a61_1[1], a61_1[0], gnd, gnd, gnd, gnd, a61_0[7], a61_0[6], a61_0[5], a61_0[4], a61_0[3], a61_0[2], a61_0[1], a61_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y61),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y61_0 = _y61[7:0];
    assign y61_1 = _y61[19:12];
    assign y61_2 = _y61[31:24];
    assign y61_3 = _y61[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y62 (
        .A({gnd, gnd, gnd, gnd, b62_3[7], b62_3[6], b62_3[5], b62_3[4], b62_3[3], b62_3[2], b62_3[1], b62_3[0], gnd, gnd, gnd, gnd, b62_2[7], b62_2[6], b62_2[5], b62_2[4], b62_2[3], b62_2[2], b62_2[1], b62_2[0], gnd, gnd, gnd, gnd, b62_1[7], b62_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b62_1[5], b62_1[4], b62_1[3], b62_1[2], b62_1[1], b62_1[0], gnd, gnd, gnd, gnd, b62_0[7], b62_0[6], b62_0[5], b62_0[4], b62_0[3], b62_0[2], b62_0[1], b62_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a62_3[7], a62_3[6], a62_3[5], a62_3[4], a62_3[3], a62_3[2], a62_3[1], a62_3[0], gnd, gnd, gnd, gnd, a62_2[7], a62_2[6], a62_2[5], a62_2[4], a62_2[3], a62_2[2], a62_2[1], a62_2[0], gnd, gnd, gnd, gnd, a62_1[7], a62_1[6], a62_1[5], a62_1[4], a62_1[3], a62_1[2], a62_1[1], a62_1[0], gnd, gnd, gnd, gnd, a62_0[7], a62_0[6], a62_0[5], a62_0[4], a62_0[3], a62_0[2], a62_0[1], a62_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y62),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y62_0 = _y62[7:0];
    assign y62_1 = _y62[19:12];
    assign y62_2 = _y62[31:24];
    assign y62_3 = _y62[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y63 (
        .A({gnd, gnd, gnd, gnd, b63_3[7], b63_3[6], b63_3[5], b63_3[4], b63_3[3], b63_3[2], b63_3[1], b63_3[0], gnd, gnd, gnd, gnd, b63_2[7], b63_2[6], b63_2[5], b63_2[4], b63_2[3], b63_2[2], b63_2[1], b63_2[0], gnd, gnd, gnd, gnd, b63_1[7], b63_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b63_1[5], b63_1[4], b63_1[3], b63_1[2], b63_1[1], b63_1[0], gnd, gnd, gnd, gnd, b63_0[7], b63_0[6], b63_0[5], b63_0[4], b63_0[3], b63_0[2], b63_0[1], b63_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a63_3[7], a63_3[6], a63_3[5], a63_3[4], a63_3[3], a63_3[2], a63_3[1], a63_3[0], gnd, gnd, gnd, gnd, a63_2[7], a63_2[6], a63_2[5], a63_2[4], a63_2[3], a63_2[2], a63_2[1], a63_2[0], gnd, gnd, gnd, gnd, a63_1[7], a63_1[6], a63_1[5], a63_1[4], a63_1[3], a63_1[2], a63_1[1], a63_1[0], gnd, gnd, gnd, gnd, a63_0[7], a63_0[6], a63_0[5], a63_0[4], a63_0[3], a63_0[2], a63_0[1], a63_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y63),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y63_0 = _y63[7:0];
    assign y63_1 = _y63[19:12];
    assign y63_2 = _y63[31:24];
    assign y63_3 = _y63[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y64 (
        .A({gnd, gnd, gnd, gnd, b64_3[7], b64_3[6], b64_3[5], b64_3[4], b64_3[3], b64_3[2], b64_3[1], b64_3[0], gnd, gnd, gnd, gnd, b64_2[7], b64_2[6], b64_2[5], b64_2[4], b64_2[3], b64_2[2], b64_2[1], b64_2[0], gnd, gnd, gnd, gnd, b64_1[7], b64_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b64_1[5], b64_1[4], b64_1[3], b64_1[2], b64_1[1], b64_1[0], gnd, gnd, gnd, gnd, b64_0[7], b64_0[6], b64_0[5], b64_0[4], b64_0[3], b64_0[2], b64_0[1], b64_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a64_3[7], a64_3[6], a64_3[5], a64_3[4], a64_3[3], a64_3[2], a64_3[1], a64_3[0], gnd, gnd, gnd, gnd, a64_2[7], a64_2[6], a64_2[5], a64_2[4], a64_2[3], a64_2[2], a64_2[1], a64_2[0], gnd, gnd, gnd, gnd, a64_1[7], a64_1[6], a64_1[5], a64_1[4], a64_1[3], a64_1[2], a64_1[1], a64_1[0], gnd, gnd, gnd, gnd, a64_0[7], a64_0[6], a64_0[5], a64_0[4], a64_0[3], a64_0[2], a64_0[1], a64_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y64),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y64_0 = _y64[7:0];
    assign y64_1 = _y64[19:12];
    assign y64_2 = _y64[31:24];
    assign y64_3 = _y64[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y65 (
        .A({gnd, gnd, gnd, gnd, b65_3[7], b65_3[6], b65_3[5], b65_3[4], b65_3[3], b65_3[2], b65_3[1], b65_3[0], gnd, gnd, gnd, gnd, b65_2[7], b65_2[6], b65_2[5], b65_2[4], b65_2[3], b65_2[2], b65_2[1], b65_2[0], gnd, gnd, gnd, gnd, b65_1[7], b65_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b65_1[5], b65_1[4], b65_1[3], b65_1[2], b65_1[1], b65_1[0], gnd, gnd, gnd, gnd, b65_0[7], b65_0[6], b65_0[5], b65_0[4], b65_0[3], b65_0[2], b65_0[1], b65_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a65_3[7], a65_3[6], a65_3[5], a65_3[4], a65_3[3], a65_3[2], a65_3[1], a65_3[0], gnd, gnd, gnd, gnd, a65_2[7], a65_2[6], a65_2[5], a65_2[4], a65_2[3], a65_2[2], a65_2[1], a65_2[0], gnd, gnd, gnd, gnd, a65_1[7], a65_1[6], a65_1[5], a65_1[4], a65_1[3], a65_1[2], a65_1[1], a65_1[0], gnd, gnd, gnd, gnd, a65_0[7], a65_0[6], a65_0[5], a65_0[4], a65_0[3], a65_0[2], a65_0[1], a65_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y65),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y65_0 = _y65[7:0];
    assign y65_1 = _y65[19:12];
    assign y65_2 = _y65[31:24];
    assign y65_3 = _y65[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y66 (
        .A({gnd, gnd, gnd, gnd, b66_3[7], b66_3[6], b66_3[5], b66_3[4], b66_3[3], b66_3[2], b66_3[1], b66_3[0], gnd, gnd, gnd, gnd, b66_2[7], b66_2[6], b66_2[5], b66_2[4], b66_2[3], b66_2[2], b66_2[1], b66_2[0], gnd, gnd, gnd, gnd, b66_1[7], b66_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b66_1[5], b66_1[4], b66_1[3], b66_1[2], b66_1[1], b66_1[0], gnd, gnd, gnd, gnd, b66_0[7], b66_0[6], b66_0[5], b66_0[4], b66_0[3], b66_0[2], b66_0[1], b66_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a66_3[7], a66_3[6], a66_3[5], a66_3[4], a66_3[3], a66_3[2], a66_3[1], a66_3[0], gnd, gnd, gnd, gnd, a66_2[7], a66_2[6], a66_2[5], a66_2[4], a66_2[3], a66_2[2], a66_2[1], a66_2[0], gnd, gnd, gnd, gnd, a66_1[7], a66_1[6], a66_1[5], a66_1[4], a66_1[3], a66_1[2], a66_1[1], a66_1[0], gnd, gnd, gnd, gnd, a66_0[7], a66_0[6], a66_0[5], a66_0[4], a66_0[3], a66_0[2], a66_0[1], a66_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y66),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y66_0 = _y66[7:0];
    assign y66_1 = _y66[19:12];
    assign y66_2 = _y66[31:24];
    assign y66_3 = _y66[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y67 (
        .A({gnd, gnd, gnd, gnd, b67_3[7], b67_3[6], b67_3[5], b67_3[4], b67_3[3], b67_3[2], b67_3[1], b67_3[0], gnd, gnd, gnd, gnd, b67_2[7], b67_2[6], b67_2[5], b67_2[4], b67_2[3], b67_2[2], b67_2[1], b67_2[0], gnd, gnd, gnd, gnd, b67_1[7], b67_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b67_1[5], b67_1[4], b67_1[3], b67_1[2], b67_1[1], b67_1[0], gnd, gnd, gnd, gnd, b67_0[7], b67_0[6], b67_0[5], b67_0[4], b67_0[3], b67_0[2], b67_0[1], b67_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a67_3[7], a67_3[6], a67_3[5], a67_3[4], a67_3[3], a67_3[2], a67_3[1], a67_3[0], gnd, gnd, gnd, gnd, a67_2[7], a67_2[6], a67_2[5], a67_2[4], a67_2[3], a67_2[2], a67_2[1], a67_2[0], gnd, gnd, gnd, gnd, a67_1[7], a67_1[6], a67_1[5], a67_1[4], a67_1[3], a67_1[2], a67_1[1], a67_1[0], gnd, gnd, gnd, gnd, a67_0[7], a67_0[6], a67_0[5], a67_0[4], a67_0[3], a67_0[2], a67_0[1], a67_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y67),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y67_0 = _y67[7:0];
    assign y67_1 = _y67[19:12];
    assign y67_2 = _y67[31:24];
    assign y67_3 = _y67[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y68 (
        .A({gnd, gnd, gnd, gnd, b68_3[7], b68_3[6], b68_3[5], b68_3[4], b68_3[3], b68_3[2], b68_3[1], b68_3[0], gnd, gnd, gnd, gnd, b68_2[7], b68_2[6], b68_2[5], b68_2[4], b68_2[3], b68_2[2], b68_2[1], b68_2[0], gnd, gnd, gnd, gnd, b68_1[7], b68_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b68_1[5], b68_1[4], b68_1[3], b68_1[2], b68_1[1], b68_1[0], gnd, gnd, gnd, gnd, b68_0[7], b68_0[6], b68_0[5], b68_0[4], b68_0[3], b68_0[2], b68_0[1], b68_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a68_3[7], a68_3[6], a68_3[5], a68_3[4], a68_3[3], a68_3[2], a68_3[1], a68_3[0], gnd, gnd, gnd, gnd, a68_2[7], a68_2[6], a68_2[5], a68_2[4], a68_2[3], a68_2[2], a68_2[1], a68_2[0], gnd, gnd, gnd, gnd, a68_1[7], a68_1[6], a68_1[5], a68_1[4], a68_1[3], a68_1[2], a68_1[1], a68_1[0], gnd, gnd, gnd, gnd, a68_0[7], a68_0[6], a68_0[5], a68_0[4], a68_0[3], a68_0[2], a68_0[1], a68_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y68),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y68_0 = _y68[7:0];
    assign y68_1 = _y68[19:12];
    assign y68_2 = _y68[31:24];
    assign y68_3 = _y68[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y69 (
        .A({gnd, gnd, gnd, gnd, b69_3[7], b69_3[6], b69_3[5], b69_3[4], b69_3[3], b69_3[2], b69_3[1], b69_3[0], gnd, gnd, gnd, gnd, b69_2[7], b69_2[6], b69_2[5], b69_2[4], b69_2[3], b69_2[2], b69_2[1], b69_2[0], gnd, gnd, gnd, gnd, b69_1[7], b69_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b69_1[5], b69_1[4], b69_1[3], b69_1[2], b69_1[1], b69_1[0], gnd, gnd, gnd, gnd, b69_0[7], b69_0[6], b69_0[5], b69_0[4], b69_0[3], b69_0[2], b69_0[1], b69_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a69_3[7], a69_3[6], a69_3[5], a69_3[4], a69_3[3], a69_3[2], a69_3[1], a69_3[0], gnd, gnd, gnd, gnd, a69_2[7], a69_2[6], a69_2[5], a69_2[4], a69_2[3], a69_2[2], a69_2[1], a69_2[0], gnd, gnd, gnd, gnd, a69_1[7], a69_1[6], a69_1[5], a69_1[4], a69_1[3], a69_1[2], a69_1[1], a69_1[0], gnd, gnd, gnd, gnd, a69_0[7], a69_0[6], a69_0[5], a69_0[4], a69_0[3], a69_0[2], a69_0[1], a69_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y69),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y69_0 = _y69[7:0];
    assign y69_1 = _y69[19:12];
    assign y69_2 = _y69[31:24];
    assign y69_3 = _y69[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y70 (
        .A({gnd, gnd, gnd, gnd, b70_3[7], b70_3[6], b70_3[5], b70_3[4], b70_3[3], b70_3[2], b70_3[1], b70_3[0], gnd, gnd, gnd, gnd, b70_2[7], b70_2[6], b70_2[5], b70_2[4], b70_2[3], b70_2[2], b70_2[1], b70_2[0], gnd, gnd, gnd, gnd, b70_1[7], b70_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b70_1[5], b70_1[4], b70_1[3], b70_1[2], b70_1[1], b70_1[0], gnd, gnd, gnd, gnd, b70_0[7], b70_0[6], b70_0[5], b70_0[4], b70_0[3], b70_0[2], b70_0[1], b70_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a70_3[7], a70_3[6], a70_3[5], a70_3[4], a70_3[3], a70_3[2], a70_3[1], a70_3[0], gnd, gnd, gnd, gnd, a70_2[7], a70_2[6], a70_2[5], a70_2[4], a70_2[3], a70_2[2], a70_2[1], a70_2[0], gnd, gnd, gnd, gnd, a70_1[7], a70_1[6], a70_1[5], a70_1[4], a70_1[3], a70_1[2], a70_1[1], a70_1[0], gnd, gnd, gnd, gnd, a70_0[7], a70_0[6], a70_0[5], a70_0[4], a70_0[3], a70_0[2], a70_0[1], a70_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y70),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y70_0 = _y70[7:0];
    assign y70_1 = _y70[19:12];
    assign y70_2 = _y70[31:24];
    assign y70_3 = _y70[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y71 (
        .A({gnd, gnd, gnd, gnd, b71_3[7], b71_3[6], b71_3[5], b71_3[4], b71_3[3], b71_3[2], b71_3[1], b71_3[0], gnd, gnd, gnd, gnd, b71_2[7], b71_2[6], b71_2[5], b71_2[4], b71_2[3], b71_2[2], b71_2[1], b71_2[0], gnd, gnd, gnd, gnd, b71_1[7], b71_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b71_1[5], b71_1[4], b71_1[3], b71_1[2], b71_1[1], b71_1[0], gnd, gnd, gnd, gnd, b71_0[7], b71_0[6], b71_0[5], b71_0[4], b71_0[3], b71_0[2], b71_0[1], b71_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a71_3[7], a71_3[6], a71_3[5], a71_3[4], a71_3[3], a71_3[2], a71_3[1], a71_3[0], gnd, gnd, gnd, gnd, a71_2[7], a71_2[6], a71_2[5], a71_2[4], a71_2[3], a71_2[2], a71_2[1], a71_2[0], gnd, gnd, gnd, gnd, a71_1[7], a71_1[6], a71_1[5], a71_1[4], a71_1[3], a71_1[2], a71_1[1], a71_1[0], gnd, gnd, gnd, gnd, a71_0[7], a71_0[6], a71_0[5], a71_0[4], a71_0[3], a71_0[2], a71_0[1], a71_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y71),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y71_0 = _y71[7:0];
    assign y71_1 = _y71[19:12];
    assign y71_2 = _y71[31:24];
    assign y71_3 = _y71[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y72 (
        .A({gnd, gnd, gnd, gnd, b72_3[7], b72_3[6], b72_3[5], b72_3[4], b72_3[3], b72_3[2], b72_3[1], b72_3[0], gnd, gnd, gnd, gnd, b72_2[7], b72_2[6], b72_2[5], b72_2[4], b72_2[3], b72_2[2], b72_2[1], b72_2[0], gnd, gnd, gnd, gnd, b72_1[7], b72_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b72_1[5], b72_1[4], b72_1[3], b72_1[2], b72_1[1], b72_1[0], gnd, gnd, gnd, gnd, b72_0[7], b72_0[6], b72_0[5], b72_0[4], b72_0[3], b72_0[2], b72_0[1], b72_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a72_3[7], a72_3[6], a72_3[5], a72_3[4], a72_3[3], a72_3[2], a72_3[1], a72_3[0], gnd, gnd, gnd, gnd, a72_2[7], a72_2[6], a72_2[5], a72_2[4], a72_2[3], a72_2[2], a72_2[1], a72_2[0], gnd, gnd, gnd, gnd, a72_1[7], a72_1[6], a72_1[5], a72_1[4], a72_1[3], a72_1[2], a72_1[1], a72_1[0], gnd, gnd, gnd, gnd, a72_0[7], a72_0[6], a72_0[5], a72_0[4], a72_0[3], a72_0[2], a72_0[1], a72_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y72),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y72_0 = _y72[7:0];
    assign y72_1 = _y72[19:12];
    assign y72_2 = _y72[31:24];
    assign y72_3 = _y72[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y73 (
        .A({gnd, gnd, gnd, gnd, b73_3[7], b73_3[6], b73_3[5], b73_3[4], b73_3[3], b73_3[2], b73_3[1], b73_3[0], gnd, gnd, gnd, gnd, b73_2[7], b73_2[6], b73_2[5], b73_2[4], b73_2[3], b73_2[2], b73_2[1], b73_2[0], gnd, gnd, gnd, gnd, b73_1[7], b73_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b73_1[5], b73_1[4], b73_1[3], b73_1[2], b73_1[1], b73_1[0], gnd, gnd, gnd, gnd, b73_0[7], b73_0[6], b73_0[5], b73_0[4], b73_0[3], b73_0[2], b73_0[1], b73_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a73_3[7], a73_3[6], a73_3[5], a73_3[4], a73_3[3], a73_3[2], a73_3[1], a73_3[0], gnd, gnd, gnd, gnd, a73_2[7], a73_2[6], a73_2[5], a73_2[4], a73_2[3], a73_2[2], a73_2[1], a73_2[0], gnd, gnd, gnd, gnd, a73_1[7], a73_1[6], a73_1[5], a73_1[4], a73_1[3], a73_1[2], a73_1[1], a73_1[0], gnd, gnd, gnd, gnd, a73_0[7], a73_0[6], a73_0[5], a73_0[4], a73_0[3], a73_0[2], a73_0[1], a73_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y73),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y73_0 = _y73[7:0];
    assign y73_1 = _y73[19:12];
    assign y73_2 = _y73[31:24];
    assign y73_3 = _y73[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y74 (
        .A({gnd, gnd, gnd, gnd, b74_3[7], b74_3[6], b74_3[5], b74_3[4], b74_3[3], b74_3[2], b74_3[1], b74_3[0], gnd, gnd, gnd, gnd, b74_2[7], b74_2[6], b74_2[5], b74_2[4], b74_2[3], b74_2[2], b74_2[1], b74_2[0], gnd, gnd, gnd, gnd, b74_1[7], b74_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b74_1[5], b74_1[4], b74_1[3], b74_1[2], b74_1[1], b74_1[0], gnd, gnd, gnd, gnd, b74_0[7], b74_0[6], b74_0[5], b74_0[4], b74_0[3], b74_0[2], b74_0[1], b74_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a74_3[7], a74_3[6], a74_3[5], a74_3[4], a74_3[3], a74_3[2], a74_3[1], a74_3[0], gnd, gnd, gnd, gnd, a74_2[7], a74_2[6], a74_2[5], a74_2[4], a74_2[3], a74_2[2], a74_2[1], a74_2[0], gnd, gnd, gnd, gnd, a74_1[7], a74_1[6], a74_1[5], a74_1[4], a74_1[3], a74_1[2], a74_1[1], a74_1[0], gnd, gnd, gnd, gnd, a74_0[7], a74_0[6], a74_0[5], a74_0[4], a74_0[3], a74_0[2], a74_0[1], a74_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y74),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y74_0 = _y74[7:0];
    assign y74_1 = _y74[19:12];
    assign y74_2 = _y74[31:24];
    assign y74_3 = _y74[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y75 (
        .A({gnd, gnd, gnd, gnd, b75_3[7], b75_3[6], b75_3[5], b75_3[4], b75_3[3], b75_3[2], b75_3[1], b75_3[0], gnd, gnd, gnd, gnd, b75_2[7], b75_2[6], b75_2[5], b75_2[4], b75_2[3], b75_2[2], b75_2[1], b75_2[0], gnd, gnd, gnd, gnd, b75_1[7], b75_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b75_1[5], b75_1[4], b75_1[3], b75_1[2], b75_1[1], b75_1[0], gnd, gnd, gnd, gnd, b75_0[7], b75_0[6], b75_0[5], b75_0[4], b75_0[3], b75_0[2], b75_0[1], b75_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a75_3[7], a75_3[6], a75_3[5], a75_3[4], a75_3[3], a75_3[2], a75_3[1], a75_3[0], gnd, gnd, gnd, gnd, a75_2[7], a75_2[6], a75_2[5], a75_2[4], a75_2[3], a75_2[2], a75_2[1], a75_2[0], gnd, gnd, gnd, gnd, a75_1[7], a75_1[6], a75_1[5], a75_1[4], a75_1[3], a75_1[2], a75_1[1], a75_1[0], gnd, gnd, gnd, gnd, a75_0[7], a75_0[6], a75_0[5], a75_0[4], a75_0[3], a75_0[2], a75_0[1], a75_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y75),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y75_0 = _y75[7:0];
    assign y75_1 = _y75[19:12];
    assign y75_2 = _y75[31:24];
    assign y75_3 = _y75[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y76 (
        .A({gnd, gnd, gnd, gnd, b76_3[7], b76_3[6], b76_3[5], b76_3[4], b76_3[3], b76_3[2], b76_3[1], b76_3[0], gnd, gnd, gnd, gnd, b76_2[7], b76_2[6], b76_2[5], b76_2[4], b76_2[3], b76_2[2], b76_2[1], b76_2[0], gnd, gnd, gnd, gnd, b76_1[7], b76_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b76_1[5], b76_1[4], b76_1[3], b76_1[2], b76_1[1], b76_1[0], gnd, gnd, gnd, gnd, b76_0[7], b76_0[6], b76_0[5], b76_0[4], b76_0[3], b76_0[2], b76_0[1], b76_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a76_3[7], a76_3[6], a76_3[5], a76_3[4], a76_3[3], a76_3[2], a76_3[1], a76_3[0], gnd, gnd, gnd, gnd, a76_2[7], a76_2[6], a76_2[5], a76_2[4], a76_2[3], a76_2[2], a76_2[1], a76_2[0], gnd, gnd, gnd, gnd, a76_1[7], a76_1[6], a76_1[5], a76_1[4], a76_1[3], a76_1[2], a76_1[1], a76_1[0], gnd, gnd, gnd, gnd, a76_0[7], a76_0[6], a76_0[5], a76_0[4], a76_0[3], a76_0[2], a76_0[1], a76_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y76),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y76_0 = _y76[7:0];
    assign y76_1 = _y76[19:12];
    assign y76_2 = _y76[31:24];
    assign y76_3 = _y76[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y77 (
        .A({gnd, gnd, gnd, gnd, b77_3[7], b77_3[6], b77_3[5], b77_3[4], b77_3[3], b77_3[2], b77_3[1], b77_3[0], gnd, gnd, gnd, gnd, b77_2[7], b77_2[6], b77_2[5], b77_2[4], b77_2[3], b77_2[2], b77_2[1], b77_2[0], gnd, gnd, gnd, gnd, b77_1[7], b77_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b77_1[5], b77_1[4], b77_1[3], b77_1[2], b77_1[1], b77_1[0], gnd, gnd, gnd, gnd, b77_0[7], b77_0[6], b77_0[5], b77_0[4], b77_0[3], b77_0[2], b77_0[1], b77_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a77_3[7], a77_3[6], a77_3[5], a77_3[4], a77_3[3], a77_3[2], a77_3[1], a77_3[0], gnd, gnd, gnd, gnd, a77_2[7], a77_2[6], a77_2[5], a77_2[4], a77_2[3], a77_2[2], a77_2[1], a77_2[0], gnd, gnd, gnd, gnd, a77_1[7], a77_1[6], a77_1[5], a77_1[4], a77_1[3], a77_1[2], a77_1[1], a77_1[0], gnd, gnd, gnd, gnd, a77_0[7], a77_0[6], a77_0[5], a77_0[4], a77_0[3], a77_0[2], a77_0[1], a77_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y77),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y77_0 = _y77[7:0];
    assign y77_1 = _y77[19:12];
    assign y77_2 = _y77[31:24];
    assign y77_3 = _y77[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y78 (
        .A({gnd, gnd, gnd, gnd, b78_3[7], b78_3[6], b78_3[5], b78_3[4], b78_3[3], b78_3[2], b78_3[1], b78_3[0], gnd, gnd, gnd, gnd, b78_2[7], b78_2[6], b78_2[5], b78_2[4], b78_2[3], b78_2[2], b78_2[1], b78_2[0], gnd, gnd, gnd, gnd, b78_1[7], b78_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b78_1[5], b78_1[4], b78_1[3], b78_1[2], b78_1[1], b78_1[0], gnd, gnd, gnd, gnd, b78_0[7], b78_0[6], b78_0[5], b78_0[4], b78_0[3], b78_0[2], b78_0[1], b78_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a78_3[7], a78_3[6], a78_3[5], a78_3[4], a78_3[3], a78_3[2], a78_3[1], a78_3[0], gnd, gnd, gnd, gnd, a78_2[7], a78_2[6], a78_2[5], a78_2[4], a78_2[3], a78_2[2], a78_2[1], a78_2[0], gnd, gnd, gnd, gnd, a78_1[7], a78_1[6], a78_1[5], a78_1[4], a78_1[3], a78_1[2], a78_1[1], a78_1[0], gnd, gnd, gnd, gnd, a78_0[7], a78_0[6], a78_0[5], a78_0[4], a78_0[3], a78_0[2], a78_0[1], a78_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y78),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y78_0 = _y78[7:0];
    assign y78_1 = _y78[19:12];
    assign y78_2 = _y78[31:24];
    assign y78_3 = _y78[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y79 (
        .A({gnd, gnd, gnd, gnd, b79_3[7], b79_3[6], b79_3[5], b79_3[4], b79_3[3], b79_3[2], b79_3[1], b79_3[0], gnd, gnd, gnd, gnd, b79_2[7], b79_2[6], b79_2[5], b79_2[4], b79_2[3], b79_2[2], b79_2[1], b79_2[0], gnd, gnd, gnd, gnd, b79_1[7], b79_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b79_1[5], b79_1[4], b79_1[3], b79_1[2], b79_1[1], b79_1[0], gnd, gnd, gnd, gnd, b79_0[7], b79_0[6], b79_0[5], b79_0[4], b79_0[3], b79_0[2], b79_0[1], b79_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a79_3[7], a79_3[6], a79_3[5], a79_3[4], a79_3[3], a79_3[2], a79_3[1], a79_3[0], gnd, gnd, gnd, gnd, a79_2[7], a79_2[6], a79_2[5], a79_2[4], a79_2[3], a79_2[2], a79_2[1], a79_2[0], gnd, gnd, gnd, gnd, a79_1[7], a79_1[6], a79_1[5], a79_1[4], a79_1[3], a79_1[2], a79_1[1], a79_1[0], gnd, gnd, gnd, gnd, a79_0[7], a79_0[6], a79_0[5], a79_0[4], a79_0[3], a79_0[2], a79_0[1], a79_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y79),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y79_0 = _y79[7:0];
    assign y79_1 = _y79[19:12];
    assign y79_2 = _y79[31:24];
    assign y79_3 = _y79[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y80 (
        .A({gnd, gnd, gnd, gnd, b80_3[7], b80_3[6], b80_3[5], b80_3[4], b80_3[3], b80_3[2], b80_3[1], b80_3[0], gnd, gnd, gnd, gnd, b80_2[7], b80_2[6], b80_2[5], b80_2[4], b80_2[3], b80_2[2], b80_2[1], b80_2[0], gnd, gnd, gnd, gnd, b80_1[7], b80_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b80_1[5], b80_1[4], b80_1[3], b80_1[2], b80_1[1], b80_1[0], gnd, gnd, gnd, gnd, b80_0[7], b80_0[6], b80_0[5], b80_0[4], b80_0[3], b80_0[2], b80_0[1], b80_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a80_3[7], a80_3[6], a80_3[5], a80_3[4], a80_3[3], a80_3[2], a80_3[1], a80_3[0], gnd, gnd, gnd, gnd, a80_2[7], a80_2[6], a80_2[5], a80_2[4], a80_2[3], a80_2[2], a80_2[1], a80_2[0], gnd, gnd, gnd, gnd, a80_1[7], a80_1[6], a80_1[5], a80_1[4], a80_1[3], a80_1[2], a80_1[1], a80_1[0], gnd, gnd, gnd, gnd, a80_0[7], a80_0[6], a80_0[5], a80_0[4], a80_0[3], a80_0[2], a80_0[1], a80_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y80),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y80_0 = _y80[7:0];
    assign y80_1 = _y80[19:12];
    assign y80_2 = _y80[31:24];
    assign y80_3 = _y80[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y81 (
        .A({gnd, gnd, gnd, gnd, b81_3[7], b81_3[6], b81_3[5], b81_3[4], b81_3[3], b81_3[2], b81_3[1], b81_3[0], gnd, gnd, gnd, gnd, b81_2[7], b81_2[6], b81_2[5], b81_2[4], b81_2[3], b81_2[2], b81_2[1], b81_2[0], gnd, gnd, gnd, gnd, b81_1[7], b81_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b81_1[5], b81_1[4], b81_1[3], b81_1[2], b81_1[1], b81_1[0], gnd, gnd, gnd, gnd, b81_0[7], b81_0[6], b81_0[5], b81_0[4], b81_0[3], b81_0[2], b81_0[1], b81_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a81_3[7], a81_3[6], a81_3[5], a81_3[4], a81_3[3], a81_3[2], a81_3[1], a81_3[0], gnd, gnd, gnd, gnd, a81_2[7], a81_2[6], a81_2[5], a81_2[4], a81_2[3], a81_2[2], a81_2[1], a81_2[0], gnd, gnd, gnd, gnd, a81_1[7], a81_1[6], a81_1[5], a81_1[4], a81_1[3], a81_1[2], a81_1[1], a81_1[0], gnd, gnd, gnd, gnd, a81_0[7], a81_0[6], a81_0[5], a81_0[4], a81_0[3], a81_0[2], a81_0[1], a81_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y81),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y81_0 = _y81[7:0];
    assign y81_1 = _y81[19:12];
    assign y81_2 = _y81[31:24];
    assign y81_3 = _y81[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y82 (
        .A({gnd, gnd, gnd, gnd, b82_3[7], b82_3[6], b82_3[5], b82_3[4], b82_3[3], b82_3[2], b82_3[1], b82_3[0], gnd, gnd, gnd, gnd, b82_2[7], b82_2[6], b82_2[5], b82_2[4], b82_2[3], b82_2[2], b82_2[1], b82_2[0], gnd, gnd, gnd, gnd, b82_1[7], b82_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b82_1[5], b82_1[4], b82_1[3], b82_1[2], b82_1[1], b82_1[0], gnd, gnd, gnd, gnd, b82_0[7], b82_0[6], b82_0[5], b82_0[4], b82_0[3], b82_0[2], b82_0[1], b82_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a82_3[7], a82_3[6], a82_3[5], a82_3[4], a82_3[3], a82_3[2], a82_3[1], a82_3[0], gnd, gnd, gnd, gnd, a82_2[7], a82_2[6], a82_2[5], a82_2[4], a82_2[3], a82_2[2], a82_2[1], a82_2[0], gnd, gnd, gnd, gnd, a82_1[7], a82_1[6], a82_1[5], a82_1[4], a82_1[3], a82_1[2], a82_1[1], a82_1[0], gnd, gnd, gnd, gnd, a82_0[7], a82_0[6], a82_0[5], a82_0[4], a82_0[3], a82_0[2], a82_0[1], a82_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y82),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y82_0 = _y82[7:0];
    assign y82_1 = _y82[19:12];
    assign y82_2 = _y82[31:24];
    assign y82_3 = _y82[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y83 (
        .A({gnd, gnd, gnd, gnd, b83_3[7], b83_3[6], b83_3[5], b83_3[4], b83_3[3], b83_3[2], b83_3[1], b83_3[0], gnd, gnd, gnd, gnd, b83_2[7], b83_2[6], b83_2[5], b83_2[4], b83_2[3], b83_2[2], b83_2[1], b83_2[0], gnd, gnd, gnd, gnd, b83_1[7], b83_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b83_1[5], b83_1[4], b83_1[3], b83_1[2], b83_1[1], b83_1[0], gnd, gnd, gnd, gnd, b83_0[7], b83_0[6], b83_0[5], b83_0[4], b83_0[3], b83_0[2], b83_0[1], b83_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a83_3[7], a83_3[6], a83_3[5], a83_3[4], a83_3[3], a83_3[2], a83_3[1], a83_3[0], gnd, gnd, gnd, gnd, a83_2[7], a83_2[6], a83_2[5], a83_2[4], a83_2[3], a83_2[2], a83_2[1], a83_2[0], gnd, gnd, gnd, gnd, a83_1[7], a83_1[6], a83_1[5], a83_1[4], a83_1[3], a83_1[2], a83_1[1], a83_1[0], gnd, gnd, gnd, gnd, a83_0[7], a83_0[6], a83_0[5], a83_0[4], a83_0[3], a83_0[2], a83_0[1], a83_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y83),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y83_0 = _y83[7:0];
    assign y83_1 = _y83[19:12];
    assign y83_2 = _y83[31:24];
    assign y83_3 = _y83[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y84 (
        .A({gnd, gnd, gnd, gnd, b84_3[7], b84_3[6], b84_3[5], b84_3[4], b84_3[3], b84_3[2], b84_3[1], b84_3[0], gnd, gnd, gnd, gnd, b84_2[7], b84_2[6], b84_2[5], b84_2[4], b84_2[3], b84_2[2], b84_2[1], b84_2[0], gnd, gnd, gnd, gnd, b84_1[7], b84_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b84_1[5], b84_1[4], b84_1[3], b84_1[2], b84_1[1], b84_1[0], gnd, gnd, gnd, gnd, b84_0[7], b84_0[6], b84_0[5], b84_0[4], b84_0[3], b84_0[2], b84_0[1], b84_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a84_3[7], a84_3[6], a84_3[5], a84_3[4], a84_3[3], a84_3[2], a84_3[1], a84_3[0], gnd, gnd, gnd, gnd, a84_2[7], a84_2[6], a84_2[5], a84_2[4], a84_2[3], a84_2[2], a84_2[1], a84_2[0], gnd, gnd, gnd, gnd, a84_1[7], a84_1[6], a84_1[5], a84_1[4], a84_1[3], a84_1[2], a84_1[1], a84_1[0], gnd, gnd, gnd, gnd, a84_0[7], a84_0[6], a84_0[5], a84_0[4], a84_0[3], a84_0[2], a84_0[1], a84_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y84),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y84_0 = _y84[7:0];
    assign y84_1 = _y84[19:12];
    assign y84_2 = _y84[31:24];
    assign y84_3 = _y84[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y85 (
        .A({gnd, gnd, gnd, gnd, b85_3[7], b85_3[6], b85_3[5], b85_3[4], b85_3[3], b85_3[2], b85_3[1], b85_3[0], gnd, gnd, gnd, gnd, b85_2[7], b85_2[6], b85_2[5], b85_2[4], b85_2[3], b85_2[2], b85_2[1], b85_2[0], gnd, gnd, gnd, gnd, b85_1[7], b85_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b85_1[5], b85_1[4], b85_1[3], b85_1[2], b85_1[1], b85_1[0], gnd, gnd, gnd, gnd, b85_0[7], b85_0[6], b85_0[5], b85_0[4], b85_0[3], b85_0[2], b85_0[1], b85_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a85_3[7], a85_3[6], a85_3[5], a85_3[4], a85_3[3], a85_3[2], a85_3[1], a85_3[0], gnd, gnd, gnd, gnd, a85_2[7], a85_2[6], a85_2[5], a85_2[4], a85_2[3], a85_2[2], a85_2[1], a85_2[0], gnd, gnd, gnd, gnd, a85_1[7], a85_1[6], a85_1[5], a85_1[4], a85_1[3], a85_1[2], a85_1[1], a85_1[0], gnd, gnd, gnd, gnd, a85_0[7], a85_0[6], a85_0[5], a85_0[4], a85_0[3], a85_0[2], a85_0[1], a85_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y85),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y85_0 = _y85[7:0];
    assign y85_1 = _y85[19:12];
    assign y85_2 = _y85[31:24];
    assign y85_3 = _y85[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y86 (
        .A({gnd, gnd, gnd, gnd, b86_3[7], b86_3[6], b86_3[5], b86_3[4], b86_3[3], b86_3[2], b86_3[1], b86_3[0], gnd, gnd, gnd, gnd, b86_2[7], b86_2[6], b86_2[5], b86_2[4], b86_2[3], b86_2[2], b86_2[1], b86_2[0], gnd, gnd, gnd, gnd, b86_1[7], b86_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b86_1[5], b86_1[4], b86_1[3], b86_1[2], b86_1[1], b86_1[0], gnd, gnd, gnd, gnd, b86_0[7], b86_0[6], b86_0[5], b86_0[4], b86_0[3], b86_0[2], b86_0[1], b86_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a86_3[7], a86_3[6], a86_3[5], a86_3[4], a86_3[3], a86_3[2], a86_3[1], a86_3[0], gnd, gnd, gnd, gnd, a86_2[7], a86_2[6], a86_2[5], a86_2[4], a86_2[3], a86_2[2], a86_2[1], a86_2[0], gnd, gnd, gnd, gnd, a86_1[7], a86_1[6], a86_1[5], a86_1[4], a86_1[3], a86_1[2], a86_1[1], a86_1[0], gnd, gnd, gnd, gnd, a86_0[7], a86_0[6], a86_0[5], a86_0[4], a86_0[3], a86_0[2], a86_0[1], a86_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y86),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y86_0 = _y86[7:0];
    assign y86_1 = _y86[19:12];
    assign y86_2 = _y86[31:24];
    assign y86_3 = _y86[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y87 (
        .A({gnd, gnd, gnd, gnd, b87_3[7], b87_3[6], b87_3[5], b87_3[4], b87_3[3], b87_3[2], b87_3[1], b87_3[0], gnd, gnd, gnd, gnd, b87_2[7], b87_2[6], b87_2[5], b87_2[4], b87_2[3], b87_2[2], b87_2[1], b87_2[0], gnd, gnd, gnd, gnd, b87_1[7], b87_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b87_1[5], b87_1[4], b87_1[3], b87_1[2], b87_1[1], b87_1[0], gnd, gnd, gnd, gnd, b87_0[7], b87_0[6], b87_0[5], b87_0[4], b87_0[3], b87_0[2], b87_0[1], b87_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a87_3[7], a87_3[6], a87_3[5], a87_3[4], a87_3[3], a87_3[2], a87_3[1], a87_3[0], gnd, gnd, gnd, gnd, a87_2[7], a87_2[6], a87_2[5], a87_2[4], a87_2[3], a87_2[2], a87_2[1], a87_2[0], gnd, gnd, gnd, gnd, a87_1[7], a87_1[6], a87_1[5], a87_1[4], a87_1[3], a87_1[2], a87_1[1], a87_1[0], gnd, gnd, gnd, gnd, a87_0[7], a87_0[6], a87_0[5], a87_0[4], a87_0[3], a87_0[2], a87_0[1], a87_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y87),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y87_0 = _y87[7:0];
    assign y87_1 = _y87[19:12];
    assign y87_2 = _y87[31:24];
    assign y87_3 = _y87[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y88 (
        .A({gnd, gnd, gnd, gnd, b88_3[7], b88_3[6], b88_3[5], b88_3[4], b88_3[3], b88_3[2], b88_3[1], b88_3[0], gnd, gnd, gnd, gnd, b88_2[7], b88_2[6], b88_2[5], b88_2[4], b88_2[3], b88_2[2], b88_2[1], b88_2[0], gnd, gnd, gnd, gnd, b88_1[7], b88_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b88_1[5], b88_1[4], b88_1[3], b88_1[2], b88_1[1], b88_1[0], gnd, gnd, gnd, gnd, b88_0[7], b88_0[6], b88_0[5], b88_0[4], b88_0[3], b88_0[2], b88_0[1], b88_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a88_3[7], a88_3[6], a88_3[5], a88_3[4], a88_3[3], a88_3[2], a88_3[1], a88_3[0], gnd, gnd, gnd, gnd, a88_2[7], a88_2[6], a88_2[5], a88_2[4], a88_2[3], a88_2[2], a88_2[1], a88_2[0], gnd, gnd, gnd, gnd, a88_1[7], a88_1[6], a88_1[5], a88_1[4], a88_1[3], a88_1[2], a88_1[1], a88_1[0], gnd, gnd, gnd, gnd, a88_0[7], a88_0[6], a88_0[5], a88_0[4], a88_0[3], a88_0[2], a88_0[1], a88_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y88),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y88_0 = _y88[7:0];
    assign y88_1 = _y88[19:12];
    assign y88_2 = _y88[31:24];
    assign y88_3 = _y88[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y89 (
        .A({gnd, gnd, gnd, gnd, b89_3[7], b89_3[6], b89_3[5], b89_3[4], b89_3[3], b89_3[2], b89_3[1], b89_3[0], gnd, gnd, gnd, gnd, b89_2[7], b89_2[6], b89_2[5], b89_2[4], b89_2[3], b89_2[2], b89_2[1], b89_2[0], gnd, gnd, gnd, gnd, b89_1[7], b89_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b89_1[5], b89_1[4], b89_1[3], b89_1[2], b89_1[1], b89_1[0], gnd, gnd, gnd, gnd, b89_0[7], b89_0[6], b89_0[5], b89_0[4], b89_0[3], b89_0[2], b89_0[1], b89_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a89_3[7], a89_3[6], a89_3[5], a89_3[4], a89_3[3], a89_3[2], a89_3[1], a89_3[0], gnd, gnd, gnd, gnd, a89_2[7], a89_2[6], a89_2[5], a89_2[4], a89_2[3], a89_2[2], a89_2[1], a89_2[0], gnd, gnd, gnd, gnd, a89_1[7], a89_1[6], a89_1[5], a89_1[4], a89_1[3], a89_1[2], a89_1[1], a89_1[0], gnd, gnd, gnd, gnd, a89_0[7], a89_0[6], a89_0[5], a89_0[4], a89_0[3], a89_0[2], a89_0[1], a89_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y89),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y89_0 = _y89[7:0];
    assign y89_1 = _y89[19:12];
    assign y89_2 = _y89[31:24];
    assign y89_3 = _y89[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y90 (
        .A({gnd, gnd, gnd, gnd, b90_3[7], b90_3[6], b90_3[5], b90_3[4], b90_3[3], b90_3[2], b90_3[1], b90_3[0], gnd, gnd, gnd, gnd, b90_2[7], b90_2[6], b90_2[5], b90_2[4], b90_2[3], b90_2[2], b90_2[1], b90_2[0], gnd, gnd, gnd, gnd, b90_1[7], b90_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b90_1[5], b90_1[4], b90_1[3], b90_1[2], b90_1[1], b90_1[0], gnd, gnd, gnd, gnd, b90_0[7], b90_0[6], b90_0[5], b90_0[4], b90_0[3], b90_0[2], b90_0[1], b90_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a90_3[7], a90_3[6], a90_3[5], a90_3[4], a90_3[3], a90_3[2], a90_3[1], a90_3[0], gnd, gnd, gnd, gnd, a90_2[7], a90_2[6], a90_2[5], a90_2[4], a90_2[3], a90_2[2], a90_2[1], a90_2[0], gnd, gnd, gnd, gnd, a90_1[7], a90_1[6], a90_1[5], a90_1[4], a90_1[3], a90_1[2], a90_1[1], a90_1[0], gnd, gnd, gnd, gnd, a90_0[7], a90_0[6], a90_0[5], a90_0[4], a90_0[3], a90_0[2], a90_0[1], a90_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y90),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y90_0 = _y90[7:0];
    assign y90_1 = _y90[19:12];
    assign y90_2 = _y90[31:24];
    assign y90_3 = _y90[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y91 (
        .A({gnd, gnd, gnd, gnd, b91_3[7], b91_3[6], b91_3[5], b91_3[4], b91_3[3], b91_3[2], b91_3[1], b91_3[0], gnd, gnd, gnd, gnd, b91_2[7], b91_2[6], b91_2[5], b91_2[4], b91_2[3], b91_2[2], b91_2[1], b91_2[0], gnd, gnd, gnd, gnd, b91_1[7], b91_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b91_1[5], b91_1[4], b91_1[3], b91_1[2], b91_1[1], b91_1[0], gnd, gnd, gnd, gnd, b91_0[7], b91_0[6], b91_0[5], b91_0[4], b91_0[3], b91_0[2], b91_0[1], b91_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a91_3[7], a91_3[6], a91_3[5], a91_3[4], a91_3[3], a91_3[2], a91_3[1], a91_3[0], gnd, gnd, gnd, gnd, a91_2[7], a91_2[6], a91_2[5], a91_2[4], a91_2[3], a91_2[2], a91_2[1], a91_2[0], gnd, gnd, gnd, gnd, a91_1[7], a91_1[6], a91_1[5], a91_1[4], a91_1[3], a91_1[2], a91_1[1], a91_1[0], gnd, gnd, gnd, gnd, a91_0[7], a91_0[6], a91_0[5], a91_0[4], a91_0[3], a91_0[2], a91_0[1], a91_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y91),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y91_0 = _y91[7:0];
    assign y91_1 = _y91[19:12];
    assign y91_2 = _y91[31:24];
    assign y91_3 = _y91[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y92 (
        .A({gnd, gnd, gnd, gnd, b92_3[7], b92_3[6], b92_3[5], b92_3[4], b92_3[3], b92_3[2], b92_3[1], b92_3[0], gnd, gnd, gnd, gnd, b92_2[7], b92_2[6], b92_2[5], b92_2[4], b92_2[3], b92_2[2], b92_2[1], b92_2[0], gnd, gnd, gnd, gnd, b92_1[7], b92_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b92_1[5], b92_1[4], b92_1[3], b92_1[2], b92_1[1], b92_1[0], gnd, gnd, gnd, gnd, b92_0[7], b92_0[6], b92_0[5], b92_0[4], b92_0[3], b92_0[2], b92_0[1], b92_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a92_3[7], a92_3[6], a92_3[5], a92_3[4], a92_3[3], a92_3[2], a92_3[1], a92_3[0], gnd, gnd, gnd, gnd, a92_2[7], a92_2[6], a92_2[5], a92_2[4], a92_2[3], a92_2[2], a92_2[1], a92_2[0], gnd, gnd, gnd, gnd, a92_1[7], a92_1[6], a92_1[5], a92_1[4], a92_1[3], a92_1[2], a92_1[1], a92_1[0], gnd, gnd, gnd, gnd, a92_0[7], a92_0[6], a92_0[5], a92_0[4], a92_0[3], a92_0[2], a92_0[1], a92_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y92),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y92_0 = _y92[7:0];
    assign y92_1 = _y92[19:12];
    assign y92_2 = _y92[31:24];
    assign y92_3 = _y92[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y93 (
        .A({gnd, gnd, gnd, gnd, b93_3[7], b93_3[6], b93_3[5], b93_3[4], b93_3[3], b93_3[2], b93_3[1], b93_3[0], gnd, gnd, gnd, gnd, b93_2[7], b93_2[6], b93_2[5], b93_2[4], b93_2[3], b93_2[2], b93_2[1], b93_2[0], gnd, gnd, gnd, gnd, b93_1[7], b93_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b93_1[5], b93_1[4], b93_1[3], b93_1[2], b93_1[1], b93_1[0], gnd, gnd, gnd, gnd, b93_0[7], b93_0[6], b93_0[5], b93_0[4], b93_0[3], b93_0[2], b93_0[1], b93_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a93_3[7], a93_3[6], a93_3[5], a93_3[4], a93_3[3], a93_3[2], a93_3[1], a93_3[0], gnd, gnd, gnd, gnd, a93_2[7], a93_2[6], a93_2[5], a93_2[4], a93_2[3], a93_2[2], a93_2[1], a93_2[0], gnd, gnd, gnd, gnd, a93_1[7], a93_1[6], a93_1[5], a93_1[4], a93_1[3], a93_1[2], a93_1[1], a93_1[0], gnd, gnd, gnd, gnd, a93_0[7], a93_0[6], a93_0[5], a93_0[4], a93_0[3], a93_0[2], a93_0[1], a93_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y93),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y93_0 = _y93[7:0];
    assign y93_1 = _y93[19:12];
    assign y93_2 = _y93[31:24];
    assign y93_3 = _y93[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y94 (
        .A({gnd, gnd, gnd, gnd, b94_3[7], b94_3[6], b94_3[5], b94_3[4], b94_3[3], b94_3[2], b94_3[1], b94_3[0], gnd, gnd, gnd, gnd, b94_2[7], b94_2[6], b94_2[5], b94_2[4], b94_2[3], b94_2[2], b94_2[1], b94_2[0], gnd, gnd, gnd, gnd, b94_1[7], b94_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b94_1[5], b94_1[4], b94_1[3], b94_1[2], b94_1[1], b94_1[0], gnd, gnd, gnd, gnd, b94_0[7], b94_0[6], b94_0[5], b94_0[4], b94_0[3], b94_0[2], b94_0[1], b94_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a94_3[7], a94_3[6], a94_3[5], a94_3[4], a94_3[3], a94_3[2], a94_3[1], a94_3[0], gnd, gnd, gnd, gnd, a94_2[7], a94_2[6], a94_2[5], a94_2[4], a94_2[3], a94_2[2], a94_2[1], a94_2[0], gnd, gnd, gnd, gnd, a94_1[7], a94_1[6], a94_1[5], a94_1[4], a94_1[3], a94_1[2], a94_1[1], a94_1[0], gnd, gnd, gnd, gnd, a94_0[7], a94_0[6], a94_0[5], a94_0[4], a94_0[3], a94_0[2], a94_0[1], a94_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y94),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y94_0 = _y94[7:0];
    assign y94_1 = _y94[19:12];
    assign y94_2 = _y94[31:24];
    assign y94_3 = _y94[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y95 (
        .A({gnd, gnd, gnd, gnd, b95_3[7], b95_3[6], b95_3[5], b95_3[4], b95_3[3], b95_3[2], b95_3[1], b95_3[0], gnd, gnd, gnd, gnd, b95_2[7], b95_2[6], b95_2[5], b95_2[4], b95_2[3], b95_2[2], b95_2[1], b95_2[0], gnd, gnd, gnd, gnd, b95_1[7], b95_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b95_1[5], b95_1[4], b95_1[3], b95_1[2], b95_1[1], b95_1[0], gnd, gnd, gnd, gnd, b95_0[7], b95_0[6], b95_0[5], b95_0[4], b95_0[3], b95_0[2], b95_0[1], b95_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a95_3[7], a95_3[6], a95_3[5], a95_3[4], a95_3[3], a95_3[2], a95_3[1], a95_3[0], gnd, gnd, gnd, gnd, a95_2[7], a95_2[6], a95_2[5], a95_2[4], a95_2[3], a95_2[2], a95_2[1], a95_2[0], gnd, gnd, gnd, gnd, a95_1[7], a95_1[6], a95_1[5], a95_1[4], a95_1[3], a95_1[2], a95_1[1], a95_1[0], gnd, gnd, gnd, gnd, a95_0[7], a95_0[6], a95_0[5], a95_0[4], a95_0[3], a95_0[2], a95_0[1], a95_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y95),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y95_0 = _y95[7:0];
    assign y95_1 = _y95[19:12];
    assign y95_2 = _y95[31:24];
    assign y95_3 = _y95[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y96 (
        .A({gnd, gnd, gnd, gnd, b96_3[7], b96_3[6], b96_3[5], b96_3[4], b96_3[3], b96_3[2], b96_3[1], b96_3[0], gnd, gnd, gnd, gnd, b96_2[7], b96_2[6], b96_2[5], b96_2[4], b96_2[3], b96_2[2], b96_2[1], b96_2[0], gnd, gnd, gnd, gnd, b96_1[7], b96_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b96_1[5], b96_1[4], b96_1[3], b96_1[2], b96_1[1], b96_1[0], gnd, gnd, gnd, gnd, b96_0[7], b96_0[6], b96_0[5], b96_0[4], b96_0[3], b96_0[2], b96_0[1], b96_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a96_3[7], a96_3[6], a96_3[5], a96_3[4], a96_3[3], a96_3[2], a96_3[1], a96_3[0], gnd, gnd, gnd, gnd, a96_2[7], a96_2[6], a96_2[5], a96_2[4], a96_2[3], a96_2[2], a96_2[1], a96_2[0], gnd, gnd, gnd, gnd, a96_1[7], a96_1[6], a96_1[5], a96_1[4], a96_1[3], a96_1[2], a96_1[1], a96_1[0], gnd, gnd, gnd, gnd, a96_0[7], a96_0[6], a96_0[5], a96_0[4], a96_0[3], a96_0[2], a96_0[1], a96_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y96),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y96_0 = _y96[7:0];
    assign y96_1 = _y96[19:12];
    assign y96_2 = _y96[31:24];
    assign y96_3 = _y96[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y97 (
        .A({gnd, gnd, gnd, gnd, b97_3[7], b97_3[6], b97_3[5], b97_3[4], b97_3[3], b97_3[2], b97_3[1], b97_3[0], gnd, gnd, gnd, gnd, b97_2[7], b97_2[6], b97_2[5], b97_2[4], b97_2[3], b97_2[2], b97_2[1], b97_2[0], gnd, gnd, gnd, gnd, b97_1[7], b97_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b97_1[5], b97_1[4], b97_1[3], b97_1[2], b97_1[1], b97_1[0], gnd, gnd, gnd, gnd, b97_0[7], b97_0[6], b97_0[5], b97_0[4], b97_0[3], b97_0[2], b97_0[1], b97_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a97_3[7], a97_3[6], a97_3[5], a97_3[4], a97_3[3], a97_3[2], a97_3[1], a97_3[0], gnd, gnd, gnd, gnd, a97_2[7], a97_2[6], a97_2[5], a97_2[4], a97_2[3], a97_2[2], a97_2[1], a97_2[0], gnd, gnd, gnd, gnd, a97_1[7], a97_1[6], a97_1[5], a97_1[4], a97_1[3], a97_1[2], a97_1[1], a97_1[0], gnd, gnd, gnd, gnd, a97_0[7], a97_0[6], a97_0[5], a97_0[4], a97_0[3], a97_0[2], a97_0[1], a97_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y97),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y97_0 = _y97[7:0];
    assign y97_1 = _y97[19:12];
    assign y97_2 = _y97[31:24];
    assign y97_3 = _y97[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y98 (
        .A({gnd, gnd, gnd, gnd, b98_3[7], b98_3[6], b98_3[5], b98_3[4], b98_3[3], b98_3[2], b98_3[1], b98_3[0], gnd, gnd, gnd, gnd, b98_2[7], b98_2[6], b98_2[5], b98_2[4], b98_2[3], b98_2[2], b98_2[1], b98_2[0], gnd, gnd, gnd, gnd, b98_1[7], b98_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b98_1[5], b98_1[4], b98_1[3], b98_1[2], b98_1[1], b98_1[0], gnd, gnd, gnd, gnd, b98_0[7], b98_0[6], b98_0[5], b98_0[4], b98_0[3], b98_0[2], b98_0[1], b98_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a98_3[7], a98_3[6], a98_3[5], a98_3[4], a98_3[3], a98_3[2], a98_3[1], a98_3[0], gnd, gnd, gnd, gnd, a98_2[7], a98_2[6], a98_2[5], a98_2[4], a98_2[3], a98_2[2], a98_2[1], a98_2[0], gnd, gnd, gnd, gnd, a98_1[7], a98_1[6], a98_1[5], a98_1[4], a98_1[3], a98_1[2], a98_1[1], a98_1[0], gnd, gnd, gnd, gnd, a98_0[7], a98_0[6], a98_0[5], a98_0[4], a98_0[3], a98_0[2], a98_0[1], a98_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y98),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y98_0 = _y98[7:0];
    assign y98_1 = _y98[19:12];
    assign y98_2 = _y98[31:24];
    assign y98_3 = _y98[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y99 (
        .A({gnd, gnd, gnd, gnd, b99_3[7], b99_3[6], b99_3[5], b99_3[4], b99_3[3], b99_3[2], b99_3[1], b99_3[0], gnd, gnd, gnd, gnd, b99_2[7], b99_2[6], b99_2[5], b99_2[4], b99_2[3], b99_2[2], b99_2[1], b99_2[0], gnd, gnd, gnd, gnd, b99_1[7], b99_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b99_1[5], b99_1[4], b99_1[3], b99_1[2], b99_1[1], b99_1[0], gnd, gnd, gnd, gnd, b99_0[7], b99_0[6], b99_0[5], b99_0[4], b99_0[3], b99_0[2], b99_0[1], b99_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a99_3[7], a99_3[6], a99_3[5], a99_3[4], a99_3[3], a99_3[2], a99_3[1], a99_3[0], gnd, gnd, gnd, gnd, a99_2[7], a99_2[6], a99_2[5], a99_2[4], a99_2[3], a99_2[2], a99_2[1], a99_2[0], gnd, gnd, gnd, gnd, a99_1[7], a99_1[6], a99_1[5], a99_1[4], a99_1[3], a99_1[2], a99_1[1], a99_1[0], gnd, gnd, gnd, gnd, a99_0[7], a99_0[6], a99_0[5], a99_0[4], a99_0[3], a99_0[2], a99_0[1], a99_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y99),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y99_0 = _y99[7:0];
    assign y99_1 = _y99[19:12];
    assign y99_2 = _y99[31:24];
    assign y99_3 = _y99[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y100 (
        .A({gnd, gnd, gnd, gnd, b100_3[7], b100_3[6], b100_3[5], b100_3[4], b100_3[3], b100_3[2], b100_3[1], b100_3[0], gnd, gnd, gnd, gnd, b100_2[7], b100_2[6], b100_2[5], b100_2[4], b100_2[3], b100_2[2], b100_2[1], b100_2[0], gnd, gnd, gnd, gnd, b100_1[7], b100_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b100_1[5], b100_1[4], b100_1[3], b100_1[2], b100_1[1], b100_1[0], gnd, gnd, gnd, gnd, b100_0[7], b100_0[6], b100_0[5], b100_0[4], b100_0[3], b100_0[2], b100_0[1], b100_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a100_3[7], a100_3[6], a100_3[5], a100_3[4], a100_3[3], a100_3[2], a100_3[1], a100_3[0], gnd, gnd, gnd, gnd, a100_2[7], a100_2[6], a100_2[5], a100_2[4], a100_2[3], a100_2[2], a100_2[1], a100_2[0], gnd, gnd, gnd, gnd, a100_1[7], a100_1[6], a100_1[5], a100_1[4], a100_1[3], a100_1[2], a100_1[1], a100_1[0], gnd, gnd, gnd, gnd, a100_0[7], a100_0[6], a100_0[5], a100_0[4], a100_0[3], a100_0[2], a100_0[1], a100_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y100),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y100_0 = _y100[7:0];
    assign y100_1 = _y100[19:12];
    assign y100_2 = _y100[31:24];
    assign y100_3 = _y100[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y101 (
        .A({gnd, gnd, gnd, gnd, b101_3[7], b101_3[6], b101_3[5], b101_3[4], b101_3[3], b101_3[2], b101_3[1], b101_3[0], gnd, gnd, gnd, gnd, b101_2[7], b101_2[6], b101_2[5], b101_2[4], b101_2[3], b101_2[2], b101_2[1], b101_2[0], gnd, gnd, gnd, gnd, b101_1[7], b101_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b101_1[5], b101_1[4], b101_1[3], b101_1[2], b101_1[1], b101_1[0], gnd, gnd, gnd, gnd, b101_0[7], b101_0[6], b101_0[5], b101_0[4], b101_0[3], b101_0[2], b101_0[1], b101_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a101_3[7], a101_3[6], a101_3[5], a101_3[4], a101_3[3], a101_3[2], a101_3[1], a101_3[0], gnd, gnd, gnd, gnd, a101_2[7], a101_2[6], a101_2[5], a101_2[4], a101_2[3], a101_2[2], a101_2[1], a101_2[0], gnd, gnd, gnd, gnd, a101_1[7], a101_1[6], a101_1[5], a101_1[4], a101_1[3], a101_1[2], a101_1[1], a101_1[0], gnd, gnd, gnd, gnd, a101_0[7], a101_0[6], a101_0[5], a101_0[4], a101_0[3], a101_0[2], a101_0[1], a101_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y101),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y101_0 = _y101[7:0];
    assign y101_1 = _y101[19:12];
    assign y101_2 = _y101[31:24];
    assign y101_3 = _y101[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y102 (
        .A({gnd, gnd, gnd, gnd, b102_3[7], b102_3[6], b102_3[5], b102_3[4], b102_3[3], b102_3[2], b102_3[1], b102_3[0], gnd, gnd, gnd, gnd, b102_2[7], b102_2[6], b102_2[5], b102_2[4], b102_2[3], b102_2[2], b102_2[1], b102_2[0], gnd, gnd, gnd, gnd, b102_1[7], b102_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b102_1[5], b102_1[4], b102_1[3], b102_1[2], b102_1[1], b102_1[0], gnd, gnd, gnd, gnd, b102_0[7], b102_0[6], b102_0[5], b102_0[4], b102_0[3], b102_0[2], b102_0[1], b102_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a102_3[7], a102_3[6], a102_3[5], a102_3[4], a102_3[3], a102_3[2], a102_3[1], a102_3[0], gnd, gnd, gnd, gnd, a102_2[7], a102_2[6], a102_2[5], a102_2[4], a102_2[3], a102_2[2], a102_2[1], a102_2[0], gnd, gnd, gnd, gnd, a102_1[7], a102_1[6], a102_1[5], a102_1[4], a102_1[3], a102_1[2], a102_1[1], a102_1[0], gnd, gnd, gnd, gnd, a102_0[7], a102_0[6], a102_0[5], a102_0[4], a102_0[3], a102_0[2], a102_0[1], a102_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y102),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y102_0 = _y102[7:0];
    assign y102_1 = _y102[19:12];
    assign y102_2 = _y102[31:24];
    assign y102_3 = _y102[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y103 (
        .A({gnd, gnd, gnd, gnd, b103_3[7], b103_3[6], b103_3[5], b103_3[4], b103_3[3], b103_3[2], b103_3[1], b103_3[0], gnd, gnd, gnd, gnd, b103_2[7], b103_2[6], b103_2[5], b103_2[4], b103_2[3], b103_2[2], b103_2[1], b103_2[0], gnd, gnd, gnd, gnd, b103_1[7], b103_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b103_1[5], b103_1[4], b103_1[3], b103_1[2], b103_1[1], b103_1[0], gnd, gnd, gnd, gnd, b103_0[7], b103_0[6], b103_0[5], b103_0[4], b103_0[3], b103_0[2], b103_0[1], b103_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a103_3[7], a103_3[6], a103_3[5], a103_3[4], a103_3[3], a103_3[2], a103_3[1], a103_3[0], gnd, gnd, gnd, gnd, a103_2[7], a103_2[6], a103_2[5], a103_2[4], a103_2[3], a103_2[2], a103_2[1], a103_2[0], gnd, gnd, gnd, gnd, a103_1[7], a103_1[6], a103_1[5], a103_1[4], a103_1[3], a103_1[2], a103_1[1], a103_1[0], gnd, gnd, gnd, gnd, a103_0[7], a103_0[6], a103_0[5], a103_0[4], a103_0[3], a103_0[2], a103_0[1], a103_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y103),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y103_0 = _y103[7:0];
    assign y103_1 = _y103[19:12];
    assign y103_2 = _y103[31:24];
    assign y103_3 = _y103[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y104 (
        .A({gnd, gnd, gnd, gnd, b104_3[7], b104_3[6], b104_3[5], b104_3[4], b104_3[3], b104_3[2], b104_3[1], b104_3[0], gnd, gnd, gnd, gnd, b104_2[7], b104_2[6], b104_2[5], b104_2[4], b104_2[3], b104_2[2], b104_2[1], b104_2[0], gnd, gnd, gnd, gnd, b104_1[7], b104_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b104_1[5], b104_1[4], b104_1[3], b104_1[2], b104_1[1], b104_1[0], gnd, gnd, gnd, gnd, b104_0[7], b104_0[6], b104_0[5], b104_0[4], b104_0[3], b104_0[2], b104_0[1], b104_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a104_3[7], a104_3[6], a104_3[5], a104_3[4], a104_3[3], a104_3[2], a104_3[1], a104_3[0], gnd, gnd, gnd, gnd, a104_2[7], a104_2[6], a104_2[5], a104_2[4], a104_2[3], a104_2[2], a104_2[1], a104_2[0], gnd, gnd, gnd, gnd, a104_1[7], a104_1[6], a104_1[5], a104_1[4], a104_1[3], a104_1[2], a104_1[1], a104_1[0], gnd, gnd, gnd, gnd, a104_0[7], a104_0[6], a104_0[5], a104_0[4], a104_0[3], a104_0[2], a104_0[1], a104_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y104),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y104_0 = _y104[7:0];
    assign y104_1 = _y104[19:12];
    assign y104_2 = _y104[31:24];
    assign y104_3 = _y104[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y105 (
        .A({gnd, gnd, gnd, gnd, b105_3[7], b105_3[6], b105_3[5], b105_3[4], b105_3[3], b105_3[2], b105_3[1], b105_3[0], gnd, gnd, gnd, gnd, b105_2[7], b105_2[6], b105_2[5], b105_2[4], b105_2[3], b105_2[2], b105_2[1], b105_2[0], gnd, gnd, gnd, gnd, b105_1[7], b105_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b105_1[5], b105_1[4], b105_1[3], b105_1[2], b105_1[1], b105_1[0], gnd, gnd, gnd, gnd, b105_0[7], b105_0[6], b105_0[5], b105_0[4], b105_0[3], b105_0[2], b105_0[1], b105_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a105_3[7], a105_3[6], a105_3[5], a105_3[4], a105_3[3], a105_3[2], a105_3[1], a105_3[0], gnd, gnd, gnd, gnd, a105_2[7], a105_2[6], a105_2[5], a105_2[4], a105_2[3], a105_2[2], a105_2[1], a105_2[0], gnd, gnd, gnd, gnd, a105_1[7], a105_1[6], a105_1[5], a105_1[4], a105_1[3], a105_1[2], a105_1[1], a105_1[0], gnd, gnd, gnd, gnd, a105_0[7], a105_0[6], a105_0[5], a105_0[4], a105_0[3], a105_0[2], a105_0[1], a105_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y105),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y105_0 = _y105[7:0];
    assign y105_1 = _y105[19:12];
    assign y105_2 = _y105[31:24];
    assign y105_3 = _y105[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y106 (
        .A({gnd, gnd, gnd, gnd, b106_3[7], b106_3[6], b106_3[5], b106_3[4], b106_3[3], b106_3[2], b106_3[1], b106_3[0], gnd, gnd, gnd, gnd, b106_2[7], b106_2[6], b106_2[5], b106_2[4], b106_2[3], b106_2[2], b106_2[1], b106_2[0], gnd, gnd, gnd, gnd, b106_1[7], b106_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b106_1[5], b106_1[4], b106_1[3], b106_1[2], b106_1[1], b106_1[0], gnd, gnd, gnd, gnd, b106_0[7], b106_0[6], b106_0[5], b106_0[4], b106_0[3], b106_0[2], b106_0[1], b106_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a106_3[7], a106_3[6], a106_3[5], a106_3[4], a106_3[3], a106_3[2], a106_3[1], a106_3[0], gnd, gnd, gnd, gnd, a106_2[7], a106_2[6], a106_2[5], a106_2[4], a106_2[3], a106_2[2], a106_2[1], a106_2[0], gnd, gnd, gnd, gnd, a106_1[7], a106_1[6], a106_1[5], a106_1[4], a106_1[3], a106_1[2], a106_1[1], a106_1[0], gnd, gnd, gnd, gnd, a106_0[7], a106_0[6], a106_0[5], a106_0[4], a106_0[3], a106_0[2], a106_0[1], a106_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y106),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y106_0 = _y106[7:0];
    assign y106_1 = _y106[19:12];
    assign y106_2 = _y106[31:24];
    assign y106_3 = _y106[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y107 (
        .A({gnd, gnd, gnd, gnd, b107_3[7], b107_3[6], b107_3[5], b107_3[4], b107_3[3], b107_3[2], b107_3[1], b107_3[0], gnd, gnd, gnd, gnd, b107_2[7], b107_2[6], b107_2[5], b107_2[4], b107_2[3], b107_2[2], b107_2[1], b107_2[0], gnd, gnd, gnd, gnd, b107_1[7], b107_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b107_1[5], b107_1[4], b107_1[3], b107_1[2], b107_1[1], b107_1[0], gnd, gnd, gnd, gnd, b107_0[7], b107_0[6], b107_0[5], b107_0[4], b107_0[3], b107_0[2], b107_0[1], b107_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a107_3[7], a107_3[6], a107_3[5], a107_3[4], a107_3[3], a107_3[2], a107_3[1], a107_3[0], gnd, gnd, gnd, gnd, a107_2[7], a107_2[6], a107_2[5], a107_2[4], a107_2[3], a107_2[2], a107_2[1], a107_2[0], gnd, gnd, gnd, gnd, a107_1[7], a107_1[6], a107_1[5], a107_1[4], a107_1[3], a107_1[2], a107_1[1], a107_1[0], gnd, gnd, gnd, gnd, a107_0[7], a107_0[6], a107_0[5], a107_0[4], a107_0[3], a107_0[2], a107_0[1], a107_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y107),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y107_0 = _y107[7:0];
    assign y107_1 = _y107[19:12];
    assign y107_2 = _y107[31:24];
    assign y107_3 = _y107[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y108 (
        .A({gnd, gnd, gnd, gnd, b108_3[7], b108_3[6], b108_3[5], b108_3[4], b108_3[3], b108_3[2], b108_3[1], b108_3[0], gnd, gnd, gnd, gnd, b108_2[7], b108_2[6], b108_2[5], b108_2[4], b108_2[3], b108_2[2], b108_2[1], b108_2[0], gnd, gnd, gnd, gnd, b108_1[7], b108_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b108_1[5], b108_1[4], b108_1[3], b108_1[2], b108_1[1], b108_1[0], gnd, gnd, gnd, gnd, b108_0[7], b108_0[6], b108_0[5], b108_0[4], b108_0[3], b108_0[2], b108_0[1], b108_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a108_3[7], a108_3[6], a108_3[5], a108_3[4], a108_3[3], a108_3[2], a108_3[1], a108_3[0], gnd, gnd, gnd, gnd, a108_2[7], a108_2[6], a108_2[5], a108_2[4], a108_2[3], a108_2[2], a108_2[1], a108_2[0], gnd, gnd, gnd, gnd, a108_1[7], a108_1[6], a108_1[5], a108_1[4], a108_1[3], a108_1[2], a108_1[1], a108_1[0], gnd, gnd, gnd, gnd, a108_0[7], a108_0[6], a108_0[5], a108_0[4], a108_0[3], a108_0[2], a108_0[1], a108_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y108),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y108_0 = _y108[7:0];
    assign y108_1 = _y108[19:12];
    assign y108_2 = _y108[31:24];
    assign y108_3 = _y108[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y109 (
        .A({gnd, gnd, gnd, gnd, b109_3[7], b109_3[6], b109_3[5], b109_3[4], b109_3[3], b109_3[2], b109_3[1], b109_3[0], gnd, gnd, gnd, gnd, b109_2[7], b109_2[6], b109_2[5], b109_2[4], b109_2[3], b109_2[2], b109_2[1], b109_2[0], gnd, gnd, gnd, gnd, b109_1[7], b109_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b109_1[5], b109_1[4], b109_1[3], b109_1[2], b109_1[1], b109_1[0], gnd, gnd, gnd, gnd, b109_0[7], b109_0[6], b109_0[5], b109_0[4], b109_0[3], b109_0[2], b109_0[1], b109_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a109_3[7], a109_3[6], a109_3[5], a109_3[4], a109_3[3], a109_3[2], a109_3[1], a109_3[0], gnd, gnd, gnd, gnd, a109_2[7], a109_2[6], a109_2[5], a109_2[4], a109_2[3], a109_2[2], a109_2[1], a109_2[0], gnd, gnd, gnd, gnd, a109_1[7], a109_1[6], a109_1[5], a109_1[4], a109_1[3], a109_1[2], a109_1[1], a109_1[0], gnd, gnd, gnd, gnd, a109_0[7], a109_0[6], a109_0[5], a109_0[4], a109_0[3], a109_0[2], a109_0[1], a109_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y109),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y109_0 = _y109[7:0];
    assign y109_1 = _y109[19:12];
    assign y109_2 = _y109[31:24];
    assign y109_3 = _y109[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y110 (
        .A({gnd, gnd, gnd, gnd, b110_3[7], b110_3[6], b110_3[5], b110_3[4], b110_3[3], b110_3[2], b110_3[1], b110_3[0], gnd, gnd, gnd, gnd, b110_2[7], b110_2[6], b110_2[5], b110_2[4], b110_2[3], b110_2[2], b110_2[1], b110_2[0], gnd, gnd, gnd, gnd, b110_1[7], b110_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b110_1[5], b110_1[4], b110_1[3], b110_1[2], b110_1[1], b110_1[0], gnd, gnd, gnd, gnd, b110_0[7], b110_0[6], b110_0[5], b110_0[4], b110_0[3], b110_0[2], b110_0[1], b110_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a110_3[7], a110_3[6], a110_3[5], a110_3[4], a110_3[3], a110_3[2], a110_3[1], a110_3[0], gnd, gnd, gnd, gnd, a110_2[7], a110_2[6], a110_2[5], a110_2[4], a110_2[3], a110_2[2], a110_2[1], a110_2[0], gnd, gnd, gnd, gnd, a110_1[7], a110_1[6], a110_1[5], a110_1[4], a110_1[3], a110_1[2], a110_1[1], a110_1[0], gnd, gnd, gnd, gnd, a110_0[7], a110_0[6], a110_0[5], a110_0[4], a110_0[3], a110_0[2], a110_0[1], a110_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y110),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y110_0 = _y110[7:0];
    assign y110_1 = _y110[19:12];
    assign y110_2 = _y110[31:24];
    assign y110_3 = _y110[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y111 (
        .A({gnd, gnd, gnd, gnd, b111_3[7], b111_3[6], b111_3[5], b111_3[4], b111_3[3], b111_3[2], b111_3[1], b111_3[0], gnd, gnd, gnd, gnd, b111_2[7], b111_2[6], b111_2[5], b111_2[4], b111_2[3], b111_2[2], b111_2[1], b111_2[0], gnd, gnd, gnd, gnd, b111_1[7], b111_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b111_1[5], b111_1[4], b111_1[3], b111_1[2], b111_1[1], b111_1[0], gnd, gnd, gnd, gnd, b111_0[7], b111_0[6], b111_0[5], b111_0[4], b111_0[3], b111_0[2], b111_0[1], b111_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a111_3[7], a111_3[6], a111_3[5], a111_3[4], a111_3[3], a111_3[2], a111_3[1], a111_3[0], gnd, gnd, gnd, gnd, a111_2[7], a111_2[6], a111_2[5], a111_2[4], a111_2[3], a111_2[2], a111_2[1], a111_2[0], gnd, gnd, gnd, gnd, a111_1[7], a111_1[6], a111_1[5], a111_1[4], a111_1[3], a111_1[2], a111_1[1], a111_1[0], gnd, gnd, gnd, gnd, a111_0[7], a111_0[6], a111_0[5], a111_0[4], a111_0[3], a111_0[2], a111_0[1], a111_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y111),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y111_0 = _y111[7:0];
    assign y111_1 = _y111[19:12];
    assign y111_2 = _y111[31:24];
    assign y111_3 = _y111[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y112 (
        .A({gnd, gnd, gnd, gnd, b112_3[7], b112_3[6], b112_3[5], b112_3[4], b112_3[3], b112_3[2], b112_3[1], b112_3[0], gnd, gnd, gnd, gnd, b112_2[7], b112_2[6], b112_2[5], b112_2[4], b112_2[3], b112_2[2], b112_2[1], b112_2[0], gnd, gnd, gnd, gnd, b112_1[7], b112_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b112_1[5], b112_1[4], b112_1[3], b112_1[2], b112_1[1], b112_1[0], gnd, gnd, gnd, gnd, b112_0[7], b112_0[6], b112_0[5], b112_0[4], b112_0[3], b112_0[2], b112_0[1], b112_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a112_3[7], a112_3[6], a112_3[5], a112_3[4], a112_3[3], a112_3[2], a112_3[1], a112_3[0], gnd, gnd, gnd, gnd, a112_2[7], a112_2[6], a112_2[5], a112_2[4], a112_2[3], a112_2[2], a112_2[1], a112_2[0], gnd, gnd, gnd, gnd, a112_1[7], a112_1[6], a112_1[5], a112_1[4], a112_1[3], a112_1[2], a112_1[1], a112_1[0], gnd, gnd, gnd, gnd, a112_0[7], a112_0[6], a112_0[5], a112_0[4], a112_0[3], a112_0[2], a112_0[1], a112_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y112),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y112_0 = _y112[7:0];
    assign y112_1 = _y112[19:12];
    assign y112_2 = _y112[31:24];
    assign y112_3 = _y112[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y113 (
        .A({gnd, gnd, gnd, gnd, b113_3[7], b113_3[6], b113_3[5], b113_3[4], b113_3[3], b113_3[2], b113_3[1], b113_3[0], gnd, gnd, gnd, gnd, b113_2[7], b113_2[6], b113_2[5], b113_2[4], b113_2[3], b113_2[2], b113_2[1], b113_2[0], gnd, gnd, gnd, gnd, b113_1[7], b113_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b113_1[5], b113_1[4], b113_1[3], b113_1[2], b113_1[1], b113_1[0], gnd, gnd, gnd, gnd, b113_0[7], b113_0[6], b113_0[5], b113_0[4], b113_0[3], b113_0[2], b113_0[1], b113_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a113_3[7], a113_3[6], a113_3[5], a113_3[4], a113_3[3], a113_3[2], a113_3[1], a113_3[0], gnd, gnd, gnd, gnd, a113_2[7], a113_2[6], a113_2[5], a113_2[4], a113_2[3], a113_2[2], a113_2[1], a113_2[0], gnd, gnd, gnd, gnd, a113_1[7], a113_1[6], a113_1[5], a113_1[4], a113_1[3], a113_1[2], a113_1[1], a113_1[0], gnd, gnd, gnd, gnd, a113_0[7], a113_0[6], a113_0[5], a113_0[4], a113_0[3], a113_0[2], a113_0[1], a113_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y113),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y113_0 = _y113[7:0];
    assign y113_1 = _y113[19:12];
    assign y113_2 = _y113[31:24];
    assign y113_3 = _y113[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y114 (
        .A({gnd, gnd, gnd, gnd, b114_3[7], b114_3[6], b114_3[5], b114_3[4], b114_3[3], b114_3[2], b114_3[1], b114_3[0], gnd, gnd, gnd, gnd, b114_2[7], b114_2[6], b114_2[5], b114_2[4], b114_2[3], b114_2[2], b114_2[1], b114_2[0], gnd, gnd, gnd, gnd, b114_1[7], b114_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b114_1[5], b114_1[4], b114_1[3], b114_1[2], b114_1[1], b114_1[0], gnd, gnd, gnd, gnd, b114_0[7], b114_0[6], b114_0[5], b114_0[4], b114_0[3], b114_0[2], b114_0[1], b114_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a114_3[7], a114_3[6], a114_3[5], a114_3[4], a114_3[3], a114_3[2], a114_3[1], a114_3[0], gnd, gnd, gnd, gnd, a114_2[7], a114_2[6], a114_2[5], a114_2[4], a114_2[3], a114_2[2], a114_2[1], a114_2[0], gnd, gnd, gnd, gnd, a114_1[7], a114_1[6], a114_1[5], a114_1[4], a114_1[3], a114_1[2], a114_1[1], a114_1[0], gnd, gnd, gnd, gnd, a114_0[7], a114_0[6], a114_0[5], a114_0[4], a114_0[3], a114_0[2], a114_0[1], a114_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y114),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y114_0 = _y114[7:0];
    assign y114_1 = _y114[19:12];
    assign y114_2 = _y114[31:24];
    assign y114_3 = _y114[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y115 (
        .A({gnd, gnd, gnd, gnd, b115_3[7], b115_3[6], b115_3[5], b115_3[4], b115_3[3], b115_3[2], b115_3[1], b115_3[0], gnd, gnd, gnd, gnd, b115_2[7], b115_2[6], b115_2[5], b115_2[4], b115_2[3], b115_2[2], b115_2[1], b115_2[0], gnd, gnd, gnd, gnd, b115_1[7], b115_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b115_1[5], b115_1[4], b115_1[3], b115_1[2], b115_1[1], b115_1[0], gnd, gnd, gnd, gnd, b115_0[7], b115_0[6], b115_0[5], b115_0[4], b115_0[3], b115_0[2], b115_0[1], b115_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a115_3[7], a115_3[6], a115_3[5], a115_3[4], a115_3[3], a115_3[2], a115_3[1], a115_3[0], gnd, gnd, gnd, gnd, a115_2[7], a115_2[6], a115_2[5], a115_2[4], a115_2[3], a115_2[2], a115_2[1], a115_2[0], gnd, gnd, gnd, gnd, a115_1[7], a115_1[6], a115_1[5], a115_1[4], a115_1[3], a115_1[2], a115_1[1], a115_1[0], gnd, gnd, gnd, gnd, a115_0[7], a115_0[6], a115_0[5], a115_0[4], a115_0[3], a115_0[2], a115_0[1], a115_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y115),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y115_0 = _y115[7:0];
    assign y115_1 = _y115[19:12];
    assign y115_2 = _y115[31:24];
    assign y115_3 = _y115[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y116 (
        .A({gnd, gnd, gnd, gnd, b116_3[7], b116_3[6], b116_3[5], b116_3[4], b116_3[3], b116_3[2], b116_3[1], b116_3[0], gnd, gnd, gnd, gnd, b116_2[7], b116_2[6], b116_2[5], b116_2[4], b116_2[3], b116_2[2], b116_2[1], b116_2[0], gnd, gnd, gnd, gnd, b116_1[7], b116_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b116_1[5], b116_1[4], b116_1[3], b116_1[2], b116_1[1], b116_1[0], gnd, gnd, gnd, gnd, b116_0[7], b116_0[6], b116_0[5], b116_0[4], b116_0[3], b116_0[2], b116_0[1], b116_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a116_3[7], a116_3[6], a116_3[5], a116_3[4], a116_3[3], a116_3[2], a116_3[1], a116_3[0], gnd, gnd, gnd, gnd, a116_2[7], a116_2[6], a116_2[5], a116_2[4], a116_2[3], a116_2[2], a116_2[1], a116_2[0], gnd, gnd, gnd, gnd, a116_1[7], a116_1[6], a116_1[5], a116_1[4], a116_1[3], a116_1[2], a116_1[1], a116_1[0], gnd, gnd, gnd, gnd, a116_0[7], a116_0[6], a116_0[5], a116_0[4], a116_0[3], a116_0[2], a116_0[1], a116_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y116),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y116_0 = _y116[7:0];
    assign y116_1 = _y116[19:12];
    assign y116_2 = _y116[31:24];
    assign y116_3 = _y116[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y117 (
        .A({gnd, gnd, gnd, gnd, b117_3[7], b117_3[6], b117_3[5], b117_3[4], b117_3[3], b117_3[2], b117_3[1], b117_3[0], gnd, gnd, gnd, gnd, b117_2[7], b117_2[6], b117_2[5], b117_2[4], b117_2[3], b117_2[2], b117_2[1], b117_2[0], gnd, gnd, gnd, gnd, b117_1[7], b117_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b117_1[5], b117_1[4], b117_1[3], b117_1[2], b117_1[1], b117_1[0], gnd, gnd, gnd, gnd, b117_0[7], b117_0[6], b117_0[5], b117_0[4], b117_0[3], b117_0[2], b117_0[1], b117_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a117_3[7], a117_3[6], a117_3[5], a117_3[4], a117_3[3], a117_3[2], a117_3[1], a117_3[0], gnd, gnd, gnd, gnd, a117_2[7], a117_2[6], a117_2[5], a117_2[4], a117_2[3], a117_2[2], a117_2[1], a117_2[0], gnd, gnd, gnd, gnd, a117_1[7], a117_1[6], a117_1[5], a117_1[4], a117_1[3], a117_1[2], a117_1[1], a117_1[0], gnd, gnd, gnd, gnd, a117_0[7], a117_0[6], a117_0[5], a117_0[4], a117_0[3], a117_0[2], a117_0[1], a117_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y117),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y117_0 = _y117[7:0];
    assign y117_1 = _y117[19:12];
    assign y117_2 = _y117[31:24];
    assign y117_3 = _y117[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y118 (
        .A({gnd, gnd, gnd, gnd, b118_3[7], b118_3[6], b118_3[5], b118_3[4], b118_3[3], b118_3[2], b118_3[1], b118_3[0], gnd, gnd, gnd, gnd, b118_2[7], b118_2[6], b118_2[5], b118_2[4], b118_2[3], b118_2[2], b118_2[1], b118_2[0], gnd, gnd, gnd, gnd, b118_1[7], b118_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b118_1[5], b118_1[4], b118_1[3], b118_1[2], b118_1[1], b118_1[0], gnd, gnd, gnd, gnd, b118_0[7], b118_0[6], b118_0[5], b118_0[4], b118_0[3], b118_0[2], b118_0[1], b118_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a118_3[7], a118_3[6], a118_3[5], a118_3[4], a118_3[3], a118_3[2], a118_3[1], a118_3[0], gnd, gnd, gnd, gnd, a118_2[7], a118_2[6], a118_2[5], a118_2[4], a118_2[3], a118_2[2], a118_2[1], a118_2[0], gnd, gnd, gnd, gnd, a118_1[7], a118_1[6], a118_1[5], a118_1[4], a118_1[3], a118_1[2], a118_1[1], a118_1[0], gnd, gnd, gnd, gnd, a118_0[7], a118_0[6], a118_0[5], a118_0[4], a118_0[3], a118_0[2], a118_0[1], a118_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y118),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y118_0 = _y118[7:0];
    assign y118_1 = _y118[19:12];
    assign y118_2 = _y118[31:24];
    assign y118_3 = _y118[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y119 (
        .A({gnd, gnd, gnd, gnd, b119_3[7], b119_3[6], b119_3[5], b119_3[4], b119_3[3], b119_3[2], b119_3[1], b119_3[0], gnd, gnd, gnd, gnd, b119_2[7], b119_2[6], b119_2[5], b119_2[4], b119_2[3], b119_2[2], b119_2[1], b119_2[0], gnd, gnd, gnd, gnd, b119_1[7], b119_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b119_1[5], b119_1[4], b119_1[3], b119_1[2], b119_1[1], b119_1[0], gnd, gnd, gnd, gnd, b119_0[7], b119_0[6], b119_0[5], b119_0[4], b119_0[3], b119_0[2], b119_0[1], b119_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a119_3[7], a119_3[6], a119_3[5], a119_3[4], a119_3[3], a119_3[2], a119_3[1], a119_3[0], gnd, gnd, gnd, gnd, a119_2[7], a119_2[6], a119_2[5], a119_2[4], a119_2[3], a119_2[2], a119_2[1], a119_2[0], gnd, gnd, gnd, gnd, a119_1[7], a119_1[6], a119_1[5], a119_1[4], a119_1[3], a119_1[2], a119_1[1], a119_1[0], gnd, gnd, gnd, gnd, a119_0[7], a119_0[6], a119_0[5], a119_0[4], a119_0[3], a119_0[2], a119_0[1], a119_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y119),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y119_0 = _y119[7:0];
    assign y119_1 = _y119[19:12];
    assign y119_2 = _y119[31:24];
    assign y119_3 = _y119[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y120 (
        .A({gnd, gnd, gnd, gnd, b120_3[7], b120_3[6], b120_3[5], b120_3[4], b120_3[3], b120_3[2], b120_3[1], b120_3[0], gnd, gnd, gnd, gnd, b120_2[7], b120_2[6], b120_2[5], b120_2[4], b120_2[3], b120_2[2], b120_2[1], b120_2[0], gnd, gnd, gnd, gnd, b120_1[7], b120_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b120_1[5], b120_1[4], b120_1[3], b120_1[2], b120_1[1], b120_1[0], gnd, gnd, gnd, gnd, b120_0[7], b120_0[6], b120_0[5], b120_0[4], b120_0[3], b120_0[2], b120_0[1], b120_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a120_3[7], a120_3[6], a120_3[5], a120_3[4], a120_3[3], a120_3[2], a120_3[1], a120_3[0], gnd, gnd, gnd, gnd, a120_2[7], a120_2[6], a120_2[5], a120_2[4], a120_2[3], a120_2[2], a120_2[1], a120_2[0], gnd, gnd, gnd, gnd, a120_1[7], a120_1[6], a120_1[5], a120_1[4], a120_1[3], a120_1[2], a120_1[1], a120_1[0], gnd, gnd, gnd, gnd, a120_0[7], a120_0[6], a120_0[5], a120_0[4], a120_0[3], a120_0[2], a120_0[1], a120_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y120),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y120_0 = _y120[7:0];
    assign y120_1 = _y120[19:12];
    assign y120_2 = _y120[31:24];
    assign y120_3 = _y120[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y121 (
        .A({gnd, gnd, gnd, gnd, b121_3[7], b121_3[6], b121_3[5], b121_3[4], b121_3[3], b121_3[2], b121_3[1], b121_3[0], gnd, gnd, gnd, gnd, b121_2[7], b121_2[6], b121_2[5], b121_2[4], b121_2[3], b121_2[2], b121_2[1], b121_2[0], gnd, gnd, gnd, gnd, b121_1[7], b121_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b121_1[5], b121_1[4], b121_1[3], b121_1[2], b121_1[1], b121_1[0], gnd, gnd, gnd, gnd, b121_0[7], b121_0[6], b121_0[5], b121_0[4], b121_0[3], b121_0[2], b121_0[1], b121_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a121_3[7], a121_3[6], a121_3[5], a121_3[4], a121_3[3], a121_3[2], a121_3[1], a121_3[0], gnd, gnd, gnd, gnd, a121_2[7], a121_2[6], a121_2[5], a121_2[4], a121_2[3], a121_2[2], a121_2[1], a121_2[0], gnd, gnd, gnd, gnd, a121_1[7], a121_1[6], a121_1[5], a121_1[4], a121_1[3], a121_1[2], a121_1[1], a121_1[0], gnd, gnd, gnd, gnd, a121_0[7], a121_0[6], a121_0[5], a121_0[4], a121_0[3], a121_0[2], a121_0[1], a121_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y121),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y121_0 = _y121[7:0];
    assign y121_1 = _y121[19:12];
    assign y121_2 = _y121[31:24];
    assign y121_3 = _y121[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y122 (
        .A({gnd, gnd, gnd, gnd, b122_3[7], b122_3[6], b122_3[5], b122_3[4], b122_3[3], b122_3[2], b122_3[1], b122_3[0], gnd, gnd, gnd, gnd, b122_2[7], b122_2[6], b122_2[5], b122_2[4], b122_2[3], b122_2[2], b122_2[1], b122_2[0], gnd, gnd, gnd, gnd, b122_1[7], b122_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b122_1[5], b122_1[4], b122_1[3], b122_1[2], b122_1[1], b122_1[0], gnd, gnd, gnd, gnd, b122_0[7], b122_0[6], b122_0[5], b122_0[4], b122_0[3], b122_0[2], b122_0[1], b122_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a122_3[7], a122_3[6], a122_3[5], a122_3[4], a122_3[3], a122_3[2], a122_3[1], a122_3[0], gnd, gnd, gnd, gnd, a122_2[7], a122_2[6], a122_2[5], a122_2[4], a122_2[3], a122_2[2], a122_2[1], a122_2[0], gnd, gnd, gnd, gnd, a122_1[7], a122_1[6], a122_1[5], a122_1[4], a122_1[3], a122_1[2], a122_1[1], a122_1[0], gnd, gnd, gnd, gnd, a122_0[7], a122_0[6], a122_0[5], a122_0[4], a122_0[3], a122_0[2], a122_0[1], a122_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y122),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y122_0 = _y122[7:0];
    assign y122_1 = _y122[19:12];
    assign y122_2 = _y122[31:24];
    assign y122_3 = _y122[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y123 (
        .A({gnd, gnd, gnd, gnd, b123_3[7], b123_3[6], b123_3[5], b123_3[4], b123_3[3], b123_3[2], b123_3[1], b123_3[0], gnd, gnd, gnd, gnd, b123_2[7], b123_2[6], b123_2[5], b123_2[4], b123_2[3], b123_2[2], b123_2[1], b123_2[0], gnd, gnd, gnd, gnd, b123_1[7], b123_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b123_1[5], b123_1[4], b123_1[3], b123_1[2], b123_1[1], b123_1[0], gnd, gnd, gnd, gnd, b123_0[7], b123_0[6], b123_0[5], b123_0[4], b123_0[3], b123_0[2], b123_0[1], b123_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a123_3[7], a123_3[6], a123_3[5], a123_3[4], a123_3[3], a123_3[2], a123_3[1], a123_3[0], gnd, gnd, gnd, gnd, a123_2[7], a123_2[6], a123_2[5], a123_2[4], a123_2[3], a123_2[2], a123_2[1], a123_2[0], gnd, gnd, gnd, gnd, a123_1[7], a123_1[6], a123_1[5], a123_1[4], a123_1[3], a123_1[2], a123_1[1], a123_1[0], gnd, gnd, gnd, gnd, a123_0[7], a123_0[6], a123_0[5], a123_0[4], a123_0[3], a123_0[2], a123_0[1], a123_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y123),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y123_0 = _y123[7:0];
    assign y123_1 = _y123[19:12];
    assign y123_2 = _y123[31:24];
    assign y123_3 = _y123[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y124 (
        .A({gnd, gnd, gnd, gnd, b124_3[7], b124_3[6], b124_3[5], b124_3[4], b124_3[3], b124_3[2], b124_3[1], b124_3[0], gnd, gnd, gnd, gnd, b124_2[7], b124_2[6], b124_2[5], b124_2[4], b124_2[3], b124_2[2], b124_2[1], b124_2[0], gnd, gnd, gnd, gnd, b124_1[7], b124_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b124_1[5], b124_1[4], b124_1[3], b124_1[2], b124_1[1], b124_1[0], gnd, gnd, gnd, gnd, b124_0[7], b124_0[6], b124_0[5], b124_0[4], b124_0[3], b124_0[2], b124_0[1], b124_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a124_3[7], a124_3[6], a124_3[5], a124_3[4], a124_3[3], a124_3[2], a124_3[1], a124_3[0], gnd, gnd, gnd, gnd, a124_2[7], a124_2[6], a124_2[5], a124_2[4], a124_2[3], a124_2[2], a124_2[1], a124_2[0], gnd, gnd, gnd, gnd, a124_1[7], a124_1[6], a124_1[5], a124_1[4], a124_1[3], a124_1[2], a124_1[1], a124_1[0], gnd, gnd, gnd, gnd, a124_0[7], a124_0[6], a124_0[5], a124_0[4], a124_0[3], a124_0[2], a124_0[1], a124_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y124),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y124_0 = _y124[7:0];
    assign y124_1 = _y124[19:12];
    assign y124_2 = _y124[31:24];
    assign y124_3 = _y124[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y125 (
        .A({gnd, gnd, gnd, gnd, b125_3[7], b125_3[6], b125_3[5], b125_3[4], b125_3[3], b125_3[2], b125_3[1], b125_3[0], gnd, gnd, gnd, gnd, b125_2[7], b125_2[6], b125_2[5], b125_2[4], b125_2[3], b125_2[2], b125_2[1], b125_2[0], gnd, gnd, gnd, gnd, b125_1[7], b125_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b125_1[5], b125_1[4], b125_1[3], b125_1[2], b125_1[1], b125_1[0], gnd, gnd, gnd, gnd, b125_0[7], b125_0[6], b125_0[5], b125_0[4], b125_0[3], b125_0[2], b125_0[1], b125_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a125_3[7], a125_3[6], a125_3[5], a125_3[4], a125_3[3], a125_3[2], a125_3[1], a125_3[0], gnd, gnd, gnd, gnd, a125_2[7], a125_2[6], a125_2[5], a125_2[4], a125_2[3], a125_2[2], a125_2[1], a125_2[0], gnd, gnd, gnd, gnd, a125_1[7], a125_1[6], a125_1[5], a125_1[4], a125_1[3], a125_1[2], a125_1[1], a125_1[0], gnd, gnd, gnd, gnd, a125_0[7], a125_0[6], a125_0[5], a125_0[4], a125_0[3], a125_0[2], a125_0[1], a125_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y125),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y125_0 = _y125[7:0];
    assign y125_1 = _y125[19:12];
    assign y125_2 = _y125[31:24];
    assign y125_3 = _y125[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y126 (
        .A({gnd, gnd, gnd, gnd, b126_3[7], b126_3[6], b126_3[5], b126_3[4], b126_3[3], b126_3[2], b126_3[1], b126_3[0], gnd, gnd, gnd, gnd, b126_2[7], b126_2[6], b126_2[5], b126_2[4], b126_2[3], b126_2[2], b126_2[1], b126_2[0], gnd, gnd, gnd, gnd, b126_1[7], b126_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b126_1[5], b126_1[4], b126_1[3], b126_1[2], b126_1[1], b126_1[0], gnd, gnd, gnd, gnd, b126_0[7], b126_0[6], b126_0[5], b126_0[4], b126_0[3], b126_0[2], b126_0[1], b126_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a126_3[7], a126_3[6], a126_3[5], a126_3[4], a126_3[3], a126_3[2], a126_3[1], a126_3[0], gnd, gnd, gnd, gnd, a126_2[7], a126_2[6], a126_2[5], a126_2[4], a126_2[3], a126_2[2], a126_2[1], a126_2[0], gnd, gnd, gnd, gnd, a126_1[7], a126_1[6], a126_1[5], a126_1[4], a126_1[3], a126_1[2], a126_1[1], a126_1[0], gnd, gnd, gnd, gnd, a126_0[7], a126_0[6], a126_0[5], a126_0[4], a126_0[3], a126_0[2], a126_0[1], a126_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y126),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y126_0 = _y126[7:0];
    assign y126_1 = _y126[19:12];
    assign y126_2 = _y126[31:24];
    assign y126_3 = _y126[43:36];
    DSP48E2 # (
        .ACASCREG(1),
        .ADREG(0),
        .ALUMODEREG(0),
        .AMULTSEL("A"),
        .AREG(1),
        .AUTORESET_PATDET("NO_RESET"),
        .AUTORESET_PRIORITY("RESET"),
        .A_INPUT("DIRECT"),
        .BCASCREG(1),
        .BMULTSEL("B"),
        .BREG(1),
        .B_INPUT("DIRECT"),
        .CARRYINREG(0),
        .CARRYINSELREG(0),
        .CREG(1),
        .DREG(0),
        .INMODEREG(0),
        .IS_ALUMODE_INVERTED(4'h0),
        .IS_CARRYIN_INVERTED(1'b0),
        .IS_CLK_INVERTED(1'b0),
        .IS_INMODE_INVERTED(5'h0),
        .IS_OPMODE_INVERTED(9'h0),
        .IS_RSTALLCARRYIN_INVERTED(1'b0),
        .IS_RSTALUMODE_INVERTED(1'b0),
        .IS_RSTA_INVERTED(1'b0),
        .IS_RSTB_INVERTED(1'b0),
        .IS_RSTCTRL_INVERTED(1'b0),
        .IS_RSTC_INVERTED(1'b0),
        .IS_RSTD_INVERTED(1'b0),
        .IS_RSTINMODE_INVERTED(1'b0),
        .IS_RSTM_INVERTED(1'b0),
        .IS_RSTP_INVERTED(1'b0),
        .MASK(48'h3fffffffffff),
        .MREG(0),
        .OPMODEREG(0),
        .PATTERN(48'h0),
        .PREADDINSEL("A"),
        .PREG(1),
        .RND(48'h0),
        .SEL_MASK("MASK"),
        .SEL_PATTERN("PATTERN"),
        .USE_MULT("NONE"),
        .USE_SIMD("FOUR12"),
        .USE_WIDEXOR("FALSE"),
        .XORSIMD("XOR24_48_96")
    ) __y127 (
        .A({gnd, gnd, gnd, gnd, b127_3[7], b127_3[6], b127_3[5], b127_3[4], b127_3[3], b127_3[2], b127_3[1], b127_3[0], gnd, gnd, gnd, gnd, b127_2[7], b127_2[6], b127_2[5], b127_2[4], b127_2[3], b127_2[2], b127_2[1], b127_2[0], gnd, gnd, gnd, gnd, b127_1[7], b127_1[6]}),
        .ACIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .ACOUT(),
        .ALUMODE({gnd, gnd, gnd, gnd}),
        .B({b127_1[5], b127_1[4], b127_1[3], b127_1[2], b127_1[1], b127_1[0], gnd, gnd, gnd, gnd, b127_0[7], b127_0[6], b127_0[5], b127_0[4], b127_0[3], b127_0[2], b127_0[1], b127_0[0]}),
        .BCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .BCOUT(),
        .C({gnd, gnd, gnd, gnd, a127_3[7], a127_3[6], a127_3[5], a127_3[4], a127_3[3], a127_3[2], a127_3[1], a127_3[0], gnd, gnd, gnd, gnd, a127_2[7], a127_2[6], a127_2[5], a127_2[4], a127_2[3], a127_2[2], a127_2[1], a127_2[0], gnd, gnd, gnd, gnd, a127_1[7], a127_1[6], a127_1[5], a127_1[4], a127_1[3], a127_1[2], a127_1[1], a127_1[0], gnd, gnd, gnd, gnd, a127_0[7], a127_0[6], a127_0[5], a127_0[4], a127_0[3], a127_0[2], a127_0[1], a127_0[0]}),
        .CARRYCASCIN(gnd),
        .CARRYCASCOUT(),
        .CARRYIN(gnd),
        .CARRYINSEL({gnd, gnd, gnd}),
        .CARRYOUT(),
        .CEA1(en),
        .CEA2(en),
        .CEAD(gnd),
        .CEALUMODE(gnd),
        .CEB1(en),
        .CEB2(en),
        .CEC(en),
        .CECARRYIN(gnd),
        .CECTRL(gnd),
        .CED(gnd),
        .CEINMODE(gnd),
        .CEM(gnd),
        .CEP(en),
        .CLK(clock),
        .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .INMODE({gnd, gnd, gnd, gnd, gnd}),
        .MULTSIGNIN(gnd),
        .MULTSIGNOUT(),
        .OPMODE({gnd, gnd, gnd, vcc, vcc, gnd, gnd, vcc, vcc}),
        .OVERFLOW(),
        .P(_y127),
        .PATTERNBDETECT(),
        .PATTERNDETECT(),
        .PCIN({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
        .PCOUT(),
        .RSTA(reset),
        .RSTALLCARRYIN(reset),
        .RSTALUMODE(reset),
        .RSTB(reset),
        .RSTC(reset),
        .RSTCTRL(reset),
        .RSTD(reset),
        .RSTINMODE(reset),
        .RSTM(reset),
        .RSTP(reset),
        .UNDERFLOW(),
        .XOROUT()
    );
    assign y127_0 = _y127[7:0];
    assign y127_1 = _y127[19:12];
    assign y127_2 = _y127[31:24];
    assign y127_3 = _y127[43:36];
endmodule
