module main (
    input wire clock,
    input wire reset,
    input wire c,
    input wire [127:0] a,
    input wire [127:0] b,
    output wire [127:0] y
);
    wire gnd;
    wire vcc;
    wire [7:0] t0;
    wire [7:0] t1;
    wire t3;
    wire t4;
    wire t5;
    wire t6;
    wire t7;
    wire t8;
    wire t9;
    wire t10;
    wire t11;
    wire t12;
    wire t13;
    wire t14;
    wire t15;
    wire t16;
    wire t17;
    wire t18;
    wire t19;
    wire t20;
    wire t21;
    wire t22;
    wire t23;
    wire t24;
    wire t25;
    wire t26;
    wire [7:0] t2;
    wire [7:0] t27;
    wire [7:0] t28;
    wire t30;
    wire t31;
    wire t32;
    wire t33;
    wire t34;
    wire t35;
    wire t36;
    wire t37;
    wire t38;
    wire t39;
    wire t40;
    wire t41;
    wire t42;
    wire t43;
    wire t44;
    wire t45;
    wire t46;
    wire t47;
    wire t48;
    wire t49;
    wire t50;
    wire t51;
    wire t52;
    wire t53;
    wire [7:0] t29;
    wire [7:0] t54;
    wire [7:0] t55;
    wire t57;
    wire t58;
    wire t59;
    wire t60;
    wire t61;
    wire t62;
    wire t63;
    wire t64;
    wire t65;
    wire t66;
    wire t67;
    wire t68;
    wire t69;
    wire t70;
    wire t71;
    wire t72;
    wire t73;
    wire t74;
    wire t75;
    wire t76;
    wire t77;
    wire t78;
    wire t79;
    wire t80;
    wire [7:0] t56;
    wire [7:0] t81;
    wire [7:0] t82;
    wire t84;
    wire t85;
    wire t86;
    wire t87;
    wire t88;
    wire t89;
    wire t90;
    wire t91;
    wire t92;
    wire t93;
    wire t94;
    wire t95;
    wire t96;
    wire t97;
    wire t98;
    wire t99;
    wire t100;
    wire t101;
    wire t102;
    wire t103;
    wire t104;
    wire t105;
    wire t106;
    wire t107;
    wire [7:0] t83;
    wire [7:0] t108;
    wire [7:0] t109;
    wire t111;
    wire t112;
    wire t113;
    wire t114;
    wire t115;
    wire t116;
    wire t117;
    wire t118;
    wire t119;
    wire t120;
    wire t121;
    wire t122;
    wire t123;
    wire t124;
    wire t125;
    wire t126;
    wire t127;
    wire t128;
    wire t129;
    wire t130;
    wire t131;
    wire t132;
    wire t133;
    wire t134;
    wire [7:0] t110;
    wire [7:0] t135;
    wire [7:0] t136;
    wire t138;
    wire t139;
    wire t140;
    wire t141;
    wire t142;
    wire t143;
    wire t144;
    wire t145;
    wire t146;
    wire t147;
    wire t148;
    wire t149;
    wire t150;
    wire t151;
    wire t152;
    wire t153;
    wire t154;
    wire t155;
    wire t156;
    wire t157;
    wire t158;
    wire t159;
    wire t160;
    wire t161;
    wire [7:0] t137;
    wire [7:0] t162;
    wire [7:0] t163;
    wire t165;
    wire t166;
    wire t167;
    wire t168;
    wire t169;
    wire t170;
    wire t171;
    wire t172;
    wire t173;
    wire t174;
    wire t175;
    wire t176;
    wire t177;
    wire t178;
    wire t179;
    wire t180;
    wire t181;
    wire t182;
    wire t183;
    wire t184;
    wire t185;
    wire t186;
    wire t187;
    wire t188;
    wire [7:0] t164;
    wire [7:0] t189;
    wire [7:0] t190;
    wire t192;
    wire t193;
    wire t194;
    wire t195;
    wire t196;
    wire t197;
    wire t198;
    wire t199;
    wire t200;
    wire t201;
    wire t202;
    wire t203;
    wire t204;
    wire t205;
    wire t206;
    wire t207;
    wire t208;
    wire t209;
    wire t210;
    wire t211;
    wire t212;
    wire t213;
    wire t214;
    wire t215;
    wire [7:0] t191;
    wire [7:0] t216;
    wire [7:0] t217;
    wire t219;
    wire t220;
    wire t221;
    wire t222;
    wire t223;
    wire t224;
    wire t225;
    wire t226;
    wire t227;
    wire t228;
    wire t229;
    wire t230;
    wire t231;
    wire t232;
    wire t233;
    wire t234;
    wire t235;
    wire t236;
    wire t237;
    wire t238;
    wire t239;
    wire t240;
    wire t241;
    wire t242;
    wire [7:0] t218;
    wire [7:0] t243;
    wire [7:0] t244;
    wire t246;
    wire t247;
    wire t248;
    wire t249;
    wire t250;
    wire t251;
    wire t252;
    wire t253;
    wire t254;
    wire t255;
    wire t256;
    wire t257;
    wire t258;
    wire t259;
    wire t260;
    wire t261;
    wire t262;
    wire t263;
    wire t264;
    wire t265;
    wire t266;
    wire t267;
    wire t268;
    wire t269;
    wire [7:0] t245;
    wire [7:0] t270;
    wire [7:0] t271;
    wire t273;
    wire t274;
    wire t275;
    wire t276;
    wire t277;
    wire t278;
    wire t279;
    wire t280;
    wire t281;
    wire t282;
    wire t283;
    wire t284;
    wire t285;
    wire t286;
    wire t287;
    wire t288;
    wire t289;
    wire t290;
    wire t291;
    wire t292;
    wire t293;
    wire t294;
    wire t295;
    wire t296;
    wire [7:0] t272;
    wire [7:0] t297;
    wire [7:0] t298;
    wire t300;
    wire t301;
    wire t302;
    wire t303;
    wire t304;
    wire t305;
    wire t306;
    wire t307;
    wire t308;
    wire t309;
    wire t310;
    wire t311;
    wire t312;
    wire t313;
    wire t314;
    wire t315;
    wire t316;
    wire t317;
    wire t318;
    wire t319;
    wire t320;
    wire t321;
    wire t322;
    wire t323;
    wire [7:0] t299;
    wire [7:0] t324;
    wire [7:0] t325;
    wire t327;
    wire t328;
    wire t329;
    wire t330;
    wire t331;
    wire t332;
    wire t333;
    wire t334;
    wire t335;
    wire t336;
    wire t337;
    wire t338;
    wire t339;
    wire t340;
    wire t341;
    wire t342;
    wire t343;
    wire t344;
    wire t345;
    wire t346;
    wire t347;
    wire t348;
    wire t349;
    wire t350;
    wire [7:0] t326;
    wire [7:0] t351;
    wire [7:0] t352;
    wire t354;
    wire t355;
    wire t356;
    wire t357;
    wire t358;
    wire t359;
    wire t360;
    wire t361;
    wire t362;
    wire t363;
    wire t364;
    wire t365;
    wire t366;
    wire t367;
    wire t368;
    wire t369;
    wire t370;
    wire t371;
    wire t372;
    wire t373;
    wire t374;
    wire t375;
    wire t376;
    wire t377;
    wire [7:0] t353;
    wire [7:0] t378;
    wire [7:0] t379;
    wire t381;
    wire t382;
    wire t383;
    wire t384;
    wire t385;
    wire t386;
    wire t387;
    wire t388;
    wire t389;
    wire t390;
    wire t391;
    wire t392;
    wire t393;
    wire t394;
    wire t395;
    wire t396;
    wire t397;
    wire t398;
    wire t399;
    wire t400;
    wire t401;
    wire t402;
    wire t403;
    wire t404;
    wire [7:0] t380;
    wire [7:0] t405;
    wire [7:0] t406;
    wire t408;
    wire t409;
    wire t410;
    wire t411;
    wire t412;
    wire t413;
    wire t414;
    wire t415;
    wire t416;
    wire t417;
    wire t418;
    wire t419;
    wire t420;
    wire t421;
    wire t422;
    wire t423;
    wire t424;
    wire t425;
    wire t426;
    wire t427;
    wire t428;
    wire t429;
    wire t430;
    wire t431;
    wire [7:0] t407;
    GND _gnd (
        .G(gnd)
    );
    VCC _vcc (
        .P(vcc)
    );
    assign t0 = a[7:0];
    assign t1 = b[7:0];
    assign t3 = t0[0];
    assign t4 = t0[1];
    assign t5 = t0[2];
    assign t6 = t0[3];
    assign t7 = t0[4];
    assign t8 = t0[5];
    assign t9 = t0[6];
    assign t10 = t0[7];
    assign t11 = t1[0];
    assign t12 = t1[1];
    assign t13 = t1[2];
    assign t14 = t1[3];
    assign t15 = t1[4];
    assign t16 = t1[5];
    assign t17 = t1[6];
    assign t18 = t1[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t19 (
        .I0(t3),
        .I1(t11),
        .I2(c),
        .O(t19)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t20 (
        .I0(t4),
        .I1(t12),
        .I2(c),
        .O(t20)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t21 (
        .I0(t5),
        .I1(t13),
        .I2(c),
        .O(t21)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t22 (
        .I0(t6),
        .I1(t14),
        .I2(c),
        .O(t22)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t23 (
        .I0(t7),
        .I1(t15),
        .I2(c),
        .O(t23)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t24 (
        .I0(t8),
        .I1(t16),
        .I2(c),
        .O(t24)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t25 (
        .I0(t9),
        .I1(t17),
        .I2(c),
        .O(t25)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t26 (
        .I0(t10),
        .I1(t18),
        .I2(c),
        .O(t26)
    );
    assign t2 = {t26, t25, t24, t23, t22, t21, t20, t19};
    assign t27 = a[15:8];
    assign t28 = b[15:8];
    assign t30 = t27[0];
    assign t31 = t27[1];
    assign t32 = t27[2];
    assign t33 = t27[3];
    assign t34 = t27[4];
    assign t35 = t27[5];
    assign t36 = t27[6];
    assign t37 = t27[7];
    assign t38 = t28[0];
    assign t39 = t28[1];
    assign t40 = t28[2];
    assign t41 = t28[3];
    assign t42 = t28[4];
    assign t43 = t28[5];
    assign t44 = t28[6];
    assign t45 = t28[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t46 (
        .I0(t30),
        .I1(t38),
        .I2(c),
        .O(t46)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t47 (
        .I0(t31),
        .I1(t39),
        .I2(c),
        .O(t47)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t48 (
        .I0(t32),
        .I1(t40),
        .I2(c),
        .O(t48)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t49 (
        .I0(t33),
        .I1(t41),
        .I2(c),
        .O(t49)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t50 (
        .I0(t34),
        .I1(t42),
        .I2(c),
        .O(t50)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t51 (
        .I0(t35),
        .I1(t43),
        .I2(c),
        .O(t51)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t52 (
        .I0(t36),
        .I1(t44),
        .I2(c),
        .O(t52)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t53 (
        .I0(t37),
        .I1(t45),
        .I2(c),
        .O(t53)
    );
    assign t29 = {t53, t52, t51, t50, t49, t48, t47, t46};
    assign t54 = a[23:16];
    assign t55 = b[23:16];
    assign t57 = t54[0];
    assign t58 = t54[1];
    assign t59 = t54[2];
    assign t60 = t54[3];
    assign t61 = t54[4];
    assign t62 = t54[5];
    assign t63 = t54[6];
    assign t64 = t54[7];
    assign t65 = t55[0];
    assign t66 = t55[1];
    assign t67 = t55[2];
    assign t68 = t55[3];
    assign t69 = t55[4];
    assign t70 = t55[5];
    assign t71 = t55[6];
    assign t72 = t55[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t73 (
        .I0(t57),
        .I1(t65),
        .I2(c),
        .O(t73)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t74 (
        .I0(t58),
        .I1(t66),
        .I2(c),
        .O(t74)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t75 (
        .I0(t59),
        .I1(t67),
        .I2(c),
        .O(t75)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t76 (
        .I0(t60),
        .I1(t68),
        .I2(c),
        .O(t76)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t77 (
        .I0(t61),
        .I1(t69),
        .I2(c),
        .O(t77)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t78 (
        .I0(t62),
        .I1(t70),
        .I2(c),
        .O(t78)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t79 (
        .I0(t63),
        .I1(t71),
        .I2(c),
        .O(t79)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t80 (
        .I0(t64),
        .I1(t72),
        .I2(c),
        .O(t80)
    );
    assign t56 = {t80, t79, t78, t77, t76, t75, t74, t73};
    assign t81 = a[31:24];
    assign t82 = b[31:24];
    assign t84 = t81[0];
    assign t85 = t81[1];
    assign t86 = t81[2];
    assign t87 = t81[3];
    assign t88 = t81[4];
    assign t89 = t81[5];
    assign t90 = t81[6];
    assign t91 = t81[7];
    assign t92 = t82[0];
    assign t93 = t82[1];
    assign t94 = t82[2];
    assign t95 = t82[3];
    assign t96 = t82[4];
    assign t97 = t82[5];
    assign t98 = t82[6];
    assign t99 = t82[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t100 (
        .I0(t84),
        .I1(t92),
        .I2(c),
        .O(t100)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t101 (
        .I0(t85),
        .I1(t93),
        .I2(c),
        .O(t101)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t102 (
        .I0(t86),
        .I1(t94),
        .I2(c),
        .O(t102)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t103 (
        .I0(t87),
        .I1(t95),
        .I2(c),
        .O(t103)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t104 (
        .I0(t88),
        .I1(t96),
        .I2(c),
        .O(t104)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t105 (
        .I0(t89),
        .I1(t97),
        .I2(c),
        .O(t105)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t106 (
        .I0(t90),
        .I1(t98),
        .I2(c),
        .O(t106)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t107 (
        .I0(t91),
        .I1(t99),
        .I2(c),
        .O(t107)
    );
    assign t83 = {t107, t106, t105, t104, t103, t102, t101, t100};
    assign t108 = a[39:32];
    assign t109 = b[39:32];
    assign t111 = t108[0];
    assign t112 = t108[1];
    assign t113 = t108[2];
    assign t114 = t108[3];
    assign t115 = t108[4];
    assign t116 = t108[5];
    assign t117 = t108[6];
    assign t118 = t108[7];
    assign t119 = t109[0];
    assign t120 = t109[1];
    assign t121 = t109[2];
    assign t122 = t109[3];
    assign t123 = t109[4];
    assign t124 = t109[5];
    assign t125 = t109[6];
    assign t126 = t109[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t127 (
        .I0(t111),
        .I1(t119),
        .I2(c),
        .O(t127)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t128 (
        .I0(t112),
        .I1(t120),
        .I2(c),
        .O(t128)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t129 (
        .I0(t113),
        .I1(t121),
        .I2(c),
        .O(t129)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t130 (
        .I0(t114),
        .I1(t122),
        .I2(c),
        .O(t130)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t131 (
        .I0(t115),
        .I1(t123),
        .I2(c),
        .O(t131)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t132 (
        .I0(t116),
        .I1(t124),
        .I2(c),
        .O(t132)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t133 (
        .I0(t117),
        .I1(t125),
        .I2(c),
        .O(t133)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t134 (
        .I0(t118),
        .I1(t126),
        .I2(c),
        .O(t134)
    );
    assign t110 = {t134, t133, t132, t131, t130, t129, t128, t127};
    assign t135 = a[47:40];
    assign t136 = b[47:40];
    assign t138 = t135[0];
    assign t139 = t135[1];
    assign t140 = t135[2];
    assign t141 = t135[3];
    assign t142 = t135[4];
    assign t143 = t135[5];
    assign t144 = t135[6];
    assign t145 = t135[7];
    assign t146 = t136[0];
    assign t147 = t136[1];
    assign t148 = t136[2];
    assign t149 = t136[3];
    assign t150 = t136[4];
    assign t151 = t136[5];
    assign t152 = t136[6];
    assign t153 = t136[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t154 (
        .I0(t138),
        .I1(t146),
        .I2(c),
        .O(t154)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t155 (
        .I0(t139),
        .I1(t147),
        .I2(c),
        .O(t155)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t156 (
        .I0(t140),
        .I1(t148),
        .I2(c),
        .O(t156)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t157 (
        .I0(t141),
        .I1(t149),
        .I2(c),
        .O(t157)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t158 (
        .I0(t142),
        .I1(t150),
        .I2(c),
        .O(t158)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t159 (
        .I0(t143),
        .I1(t151),
        .I2(c),
        .O(t159)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t160 (
        .I0(t144),
        .I1(t152),
        .I2(c),
        .O(t160)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t161 (
        .I0(t145),
        .I1(t153),
        .I2(c),
        .O(t161)
    );
    assign t137 = {t161, t160, t159, t158, t157, t156, t155, t154};
    assign t162 = a[55:48];
    assign t163 = b[55:48];
    assign t165 = t162[0];
    assign t166 = t162[1];
    assign t167 = t162[2];
    assign t168 = t162[3];
    assign t169 = t162[4];
    assign t170 = t162[5];
    assign t171 = t162[6];
    assign t172 = t162[7];
    assign t173 = t163[0];
    assign t174 = t163[1];
    assign t175 = t163[2];
    assign t176 = t163[3];
    assign t177 = t163[4];
    assign t178 = t163[5];
    assign t179 = t163[6];
    assign t180 = t163[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t181 (
        .I0(t165),
        .I1(t173),
        .I2(c),
        .O(t181)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t182 (
        .I0(t166),
        .I1(t174),
        .I2(c),
        .O(t182)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t183 (
        .I0(t167),
        .I1(t175),
        .I2(c),
        .O(t183)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t184 (
        .I0(t168),
        .I1(t176),
        .I2(c),
        .O(t184)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t185 (
        .I0(t169),
        .I1(t177),
        .I2(c),
        .O(t185)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t186 (
        .I0(t170),
        .I1(t178),
        .I2(c),
        .O(t186)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t187 (
        .I0(t171),
        .I1(t179),
        .I2(c),
        .O(t187)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t188 (
        .I0(t172),
        .I1(t180),
        .I2(c),
        .O(t188)
    );
    assign t164 = {t188, t187, t186, t185, t184, t183, t182, t181};
    assign t189 = a[63:56];
    assign t190 = b[63:56];
    assign t192 = t189[0];
    assign t193 = t189[1];
    assign t194 = t189[2];
    assign t195 = t189[3];
    assign t196 = t189[4];
    assign t197 = t189[5];
    assign t198 = t189[6];
    assign t199 = t189[7];
    assign t200 = t190[0];
    assign t201 = t190[1];
    assign t202 = t190[2];
    assign t203 = t190[3];
    assign t204 = t190[4];
    assign t205 = t190[5];
    assign t206 = t190[6];
    assign t207 = t190[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t208 (
        .I0(t192),
        .I1(t200),
        .I2(c),
        .O(t208)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t209 (
        .I0(t193),
        .I1(t201),
        .I2(c),
        .O(t209)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t210 (
        .I0(t194),
        .I1(t202),
        .I2(c),
        .O(t210)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t211 (
        .I0(t195),
        .I1(t203),
        .I2(c),
        .O(t211)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t212 (
        .I0(t196),
        .I1(t204),
        .I2(c),
        .O(t212)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t213 (
        .I0(t197),
        .I1(t205),
        .I2(c),
        .O(t213)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t214 (
        .I0(t198),
        .I1(t206),
        .I2(c),
        .O(t214)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t215 (
        .I0(t199),
        .I1(t207),
        .I2(c),
        .O(t215)
    );
    assign t191 = {t215, t214, t213, t212, t211, t210, t209, t208};
    assign t216 = a[71:64];
    assign t217 = b[71:64];
    assign t219 = t216[0];
    assign t220 = t216[1];
    assign t221 = t216[2];
    assign t222 = t216[3];
    assign t223 = t216[4];
    assign t224 = t216[5];
    assign t225 = t216[6];
    assign t226 = t216[7];
    assign t227 = t217[0];
    assign t228 = t217[1];
    assign t229 = t217[2];
    assign t230 = t217[3];
    assign t231 = t217[4];
    assign t232 = t217[5];
    assign t233 = t217[6];
    assign t234 = t217[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t235 (
        .I0(t219),
        .I1(t227),
        .I2(c),
        .O(t235)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t236 (
        .I0(t220),
        .I1(t228),
        .I2(c),
        .O(t236)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t237 (
        .I0(t221),
        .I1(t229),
        .I2(c),
        .O(t237)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t238 (
        .I0(t222),
        .I1(t230),
        .I2(c),
        .O(t238)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t239 (
        .I0(t223),
        .I1(t231),
        .I2(c),
        .O(t239)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t240 (
        .I0(t224),
        .I1(t232),
        .I2(c),
        .O(t240)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t241 (
        .I0(t225),
        .I1(t233),
        .I2(c),
        .O(t241)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t242 (
        .I0(t226),
        .I1(t234),
        .I2(c),
        .O(t242)
    );
    assign t218 = {t242, t241, t240, t239, t238, t237, t236, t235};
    assign t243 = a[79:72];
    assign t244 = b[79:72];
    assign t246 = t243[0];
    assign t247 = t243[1];
    assign t248 = t243[2];
    assign t249 = t243[3];
    assign t250 = t243[4];
    assign t251 = t243[5];
    assign t252 = t243[6];
    assign t253 = t243[7];
    assign t254 = t244[0];
    assign t255 = t244[1];
    assign t256 = t244[2];
    assign t257 = t244[3];
    assign t258 = t244[4];
    assign t259 = t244[5];
    assign t260 = t244[6];
    assign t261 = t244[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t262 (
        .I0(t246),
        .I1(t254),
        .I2(c),
        .O(t262)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t263 (
        .I0(t247),
        .I1(t255),
        .I2(c),
        .O(t263)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t264 (
        .I0(t248),
        .I1(t256),
        .I2(c),
        .O(t264)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t265 (
        .I0(t249),
        .I1(t257),
        .I2(c),
        .O(t265)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t266 (
        .I0(t250),
        .I1(t258),
        .I2(c),
        .O(t266)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t267 (
        .I0(t251),
        .I1(t259),
        .I2(c),
        .O(t267)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t268 (
        .I0(t252),
        .I1(t260),
        .I2(c),
        .O(t268)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t269 (
        .I0(t253),
        .I1(t261),
        .I2(c),
        .O(t269)
    );
    assign t245 = {t269, t268, t267, t266, t265, t264, t263, t262};
    assign t270 = a[87:80];
    assign t271 = b[87:80];
    assign t273 = t270[0];
    assign t274 = t270[1];
    assign t275 = t270[2];
    assign t276 = t270[3];
    assign t277 = t270[4];
    assign t278 = t270[5];
    assign t279 = t270[6];
    assign t280 = t270[7];
    assign t281 = t271[0];
    assign t282 = t271[1];
    assign t283 = t271[2];
    assign t284 = t271[3];
    assign t285 = t271[4];
    assign t286 = t271[5];
    assign t287 = t271[6];
    assign t288 = t271[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t289 (
        .I0(t273),
        .I1(t281),
        .I2(c),
        .O(t289)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t290 (
        .I0(t274),
        .I1(t282),
        .I2(c),
        .O(t290)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t291 (
        .I0(t275),
        .I1(t283),
        .I2(c),
        .O(t291)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t292 (
        .I0(t276),
        .I1(t284),
        .I2(c),
        .O(t292)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t293 (
        .I0(t277),
        .I1(t285),
        .I2(c),
        .O(t293)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t294 (
        .I0(t278),
        .I1(t286),
        .I2(c),
        .O(t294)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t295 (
        .I0(t279),
        .I1(t287),
        .I2(c),
        .O(t295)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t296 (
        .I0(t280),
        .I1(t288),
        .I2(c),
        .O(t296)
    );
    assign t272 = {t296, t295, t294, t293, t292, t291, t290, t289};
    assign t297 = a[95:88];
    assign t298 = b[95:88];
    assign t300 = t297[0];
    assign t301 = t297[1];
    assign t302 = t297[2];
    assign t303 = t297[3];
    assign t304 = t297[4];
    assign t305 = t297[5];
    assign t306 = t297[6];
    assign t307 = t297[7];
    assign t308 = t298[0];
    assign t309 = t298[1];
    assign t310 = t298[2];
    assign t311 = t298[3];
    assign t312 = t298[4];
    assign t313 = t298[5];
    assign t314 = t298[6];
    assign t315 = t298[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t316 (
        .I0(t300),
        .I1(t308),
        .I2(c),
        .O(t316)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t317 (
        .I0(t301),
        .I1(t309),
        .I2(c),
        .O(t317)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t318 (
        .I0(t302),
        .I1(t310),
        .I2(c),
        .O(t318)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t319 (
        .I0(t303),
        .I1(t311),
        .I2(c),
        .O(t319)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t320 (
        .I0(t304),
        .I1(t312),
        .I2(c),
        .O(t320)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t321 (
        .I0(t305),
        .I1(t313),
        .I2(c),
        .O(t321)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t322 (
        .I0(t306),
        .I1(t314),
        .I2(c),
        .O(t322)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t323 (
        .I0(t307),
        .I1(t315),
        .I2(c),
        .O(t323)
    );
    assign t299 = {t323, t322, t321, t320, t319, t318, t317, t316};
    assign t324 = a[103:96];
    assign t325 = b[103:96];
    assign t327 = t324[0];
    assign t328 = t324[1];
    assign t329 = t324[2];
    assign t330 = t324[3];
    assign t331 = t324[4];
    assign t332 = t324[5];
    assign t333 = t324[6];
    assign t334 = t324[7];
    assign t335 = t325[0];
    assign t336 = t325[1];
    assign t337 = t325[2];
    assign t338 = t325[3];
    assign t339 = t325[4];
    assign t340 = t325[5];
    assign t341 = t325[6];
    assign t342 = t325[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t343 (
        .I0(t327),
        .I1(t335),
        .I2(c),
        .O(t343)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t344 (
        .I0(t328),
        .I1(t336),
        .I2(c),
        .O(t344)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t345 (
        .I0(t329),
        .I1(t337),
        .I2(c),
        .O(t345)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t346 (
        .I0(t330),
        .I1(t338),
        .I2(c),
        .O(t346)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t347 (
        .I0(t331),
        .I1(t339),
        .I2(c),
        .O(t347)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t348 (
        .I0(t332),
        .I1(t340),
        .I2(c),
        .O(t348)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t349 (
        .I0(t333),
        .I1(t341),
        .I2(c),
        .O(t349)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t350 (
        .I0(t334),
        .I1(t342),
        .I2(c),
        .O(t350)
    );
    assign t326 = {t350, t349, t348, t347, t346, t345, t344, t343};
    assign t351 = a[111:104];
    assign t352 = b[111:104];
    assign t354 = t351[0];
    assign t355 = t351[1];
    assign t356 = t351[2];
    assign t357 = t351[3];
    assign t358 = t351[4];
    assign t359 = t351[5];
    assign t360 = t351[6];
    assign t361 = t351[7];
    assign t362 = t352[0];
    assign t363 = t352[1];
    assign t364 = t352[2];
    assign t365 = t352[3];
    assign t366 = t352[4];
    assign t367 = t352[5];
    assign t368 = t352[6];
    assign t369 = t352[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t370 (
        .I0(t354),
        .I1(t362),
        .I2(c),
        .O(t370)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t371 (
        .I0(t355),
        .I1(t363),
        .I2(c),
        .O(t371)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t372 (
        .I0(t356),
        .I1(t364),
        .I2(c),
        .O(t372)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t373 (
        .I0(t357),
        .I1(t365),
        .I2(c),
        .O(t373)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t374 (
        .I0(t358),
        .I1(t366),
        .I2(c),
        .O(t374)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t375 (
        .I0(t359),
        .I1(t367),
        .I2(c),
        .O(t375)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t376 (
        .I0(t360),
        .I1(t368),
        .I2(c),
        .O(t376)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t377 (
        .I0(t361),
        .I1(t369),
        .I2(c),
        .O(t377)
    );
    assign t353 = {t377, t376, t375, t374, t373, t372, t371, t370};
    assign t378 = a[119:112];
    assign t379 = b[119:112];
    assign t381 = t378[0];
    assign t382 = t378[1];
    assign t383 = t378[2];
    assign t384 = t378[3];
    assign t385 = t378[4];
    assign t386 = t378[5];
    assign t387 = t378[6];
    assign t388 = t378[7];
    assign t389 = t379[0];
    assign t390 = t379[1];
    assign t391 = t379[2];
    assign t392 = t379[3];
    assign t393 = t379[4];
    assign t394 = t379[5];
    assign t395 = t379[6];
    assign t396 = t379[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t397 (
        .I0(t381),
        .I1(t389),
        .I2(c),
        .O(t397)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t398 (
        .I0(t382),
        .I1(t390),
        .I2(c),
        .O(t398)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t399 (
        .I0(t383),
        .I1(t391),
        .I2(c),
        .O(t399)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t400 (
        .I0(t384),
        .I1(t392),
        .I2(c),
        .O(t400)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t401 (
        .I0(t385),
        .I1(t393),
        .I2(c),
        .O(t401)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t402 (
        .I0(t386),
        .I1(t394),
        .I2(c),
        .O(t402)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t403 (
        .I0(t387),
        .I1(t395),
        .I2(c),
        .O(t403)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t404 (
        .I0(t388),
        .I1(t396),
        .I2(c),
        .O(t404)
    );
    assign t380 = {t404, t403, t402, t401, t400, t399, t398, t397};
    assign t405 = a[127:120];
    assign t406 = b[127:120];
    assign t408 = t405[0];
    assign t409 = t405[1];
    assign t410 = t405[2];
    assign t411 = t405[3];
    assign t412 = t405[4];
    assign t413 = t405[5];
    assign t414 = t405[6];
    assign t415 = t405[7];
    assign t416 = t406[0];
    assign t417 = t406[1];
    assign t418 = t406[2];
    assign t419 = t406[3];
    assign t420 = t406[4];
    assign t421 = t406[5];
    assign t422 = t406[6];
    assign t423 = t406[7];
    LUT3 # (
        .INIT(8'hac)
    ) __t424 (
        .I0(t408),
        .I1(t416),
        .I2(c),
        .O(t424)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t425 (
        .I0(t409),
        .I1(t417),
        .I2(c),
        .O(t425)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t426 (
        .I0(t410),
        .I1(t418),
        .I2(c),
        .O(t426)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t427 (
        .I0(t411),
        .I1(t419),
        .I2(c),
        .O(t427)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t428 (
        .I0(t412),
        .I1(t420),
        .I2(c),
        .O(t428)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t429 (
        .I0(t413),
        .I1(t421),
        .I2(c),
        .O(t429)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t430 (
        .I0(t414),
        .I1(t422),
        .I2(c),
        .O(t430)
    );
    LUT3 # (
        .INIT(8'hac)
    ) __t431 (
        .I0(t415),
        .I1(t423),
        .I2(c),
        .O(t431)
    );
    assign t407 = {t431, t430, t429, t428, t427, t426, t425, t424};
    assign y = {t407, t380, t353, t326, t299, t272, t245, t218, t191, t164, t137, t110, t83, t56, t29, t2};
endmodule
